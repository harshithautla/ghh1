magic
tech scmos
timestamp 1554027465
<< rotate >>
rect 154 157 165 159
rect 421 157 432 159
rect 688 157 699 159
rect 131 153 133 155
rect 154 150 168 157
rect 398 153 400 155
rect 421 150 435 157
rect 665 153 667 155
rect 688 150 702 157
rect 157 148 168 150
rect 424 148 435 150
rect 691 148 702 150
rect 154 13 165 15
rect 421 13 432 15
rect 688 13 699 15
rect 131 9 133 11
rect 154 6 168 13
rect 398 9 400 11
rect 421 6 435 13
rect 665 9 667 11
rect 559 6 570 8
rect 688 6 702 13
rect 157 4 168 6
rect 424 4 435 6
rect 533 1 535 3
rect 556 -1 570 6
rect 691 4 702 6
rect 556 -3 567 -1
rect 559 -138 570 -136
rect 533 -143 535 -141
rect 556 -145 570 -138
rect 556 -147 567 -145
<< ab >>
rect 4 280 261 294
rect 4 276 86 280
rect 88 276 258 280
rect 260 276 261 280
rect 4 168 261 276
rect 4 164 86 168
rect 88 164 258 168
rect 260 164 261 168
rect 4 136 261 164
rect 4 132 86 136
rect 88 132 258 136
rect 260 132 261 136
rect 4 24 261 132
rect 4 20 86 24
rect 88 20 258 24
rect 260 20 261 24
rect 4 6 261 20
rect 263 286 528 294
rect 263 230 304 286
rect 309 280 528 286
rect 309 276 353 280
rect 355 276 525 280
rect 527 276 528 280
rect 309 254 528 276
rect 306 230 528 254
rect 263 214 528 230
rect 263 183 304 214
rect 306 190 528 214
rect 305 183 528 190
rect 263 180 528 183
rect 263 158 304 180
rect 305 168 528 180
rect 305 164 353 168
rect 355 164 525 168
rect 527 164 528 168
rect 305 158 528 164
rect 263 142 528 158
rect 263 86 304 142
rect 305 136 528 142
rect 305 132 353 136
rect 355 132 525 136
rect 527 132 528 136
rect 305 110 528 132
rect 309 86 528 110
rect 263 70 528 86
rect 263 39 304 70
rect 263 36 305 39
rect 263 14 304 36
rect 309 24 528 70
rect 309 20 353 24
rect 355 20 525 24
rect 527 20 528 24
rect 309 14 528 20
rect 263 6 528 14
rect 530 286 795 294
rect 530 230 571 286
rect 576 280 795 286
rect 576 276 620 280
rect 622 276 792 280
rect 794 276 795 280
rect 576 254 795 276
rect 573 230 795 254
rect 530 214 795 230
rect 530 190 571 214
rect 573 190 795 214
rect 530 168 795 190
rect 530 164 620 168
rect 622 164 792 168
rect 794 164 795 168
rect 530 136 795 164
rect 530 132 620 136
rect 622 132 792 136
rect 794 132 795 136
rect 530 110 795 132
rect 530 86 571 110
rect 573 86 795 110
rect 530 70 795 86
rect 530 39 571 70
rect 573 46 795 70
rect 530 36 572 39
rect 530 14 571 36
rect 576 24 795 46
rect 576 20 620 24
rect 622 20 792 24
rect 794 20 795 24
rect 576 14 795 20
rect 530 6 795 14
rect 797 183 838 294
rect 797 180 839 183
rect 797 39 838 180
rect 797 36 839 39
rect 797 6 838 36
rect 2 1 663 6
rect 2 -2 420 1
rect 422 -8 663 1
rect 422 -12 488 -8
rect 490 -12 660 -8
rect 662 -12 663 -8
rect 422 -48 663 -12
rect 665 -24 706 6
rect 665 -27 707 -24
rect 422 -53 664 -48
rect 422 -79 663 -53
rect 422 -84 664 -79
rect 422 -120 663 -84
rect 422 -124 488 -120
rect 490 -124 660 -120
rect 662 -124 663 -120
rect 422 -152 663 -124
rect 422 -156 488 -152
rect 490 -156 660 -152
rect 662 -156 663 -152
rect 422 -191 663 -156
rect 665 -168 706 -27
rect 708 -131 836 6
rect 708 -145 837 -131
rect 665 -171 707 -168
rect 422 -197 664 -191
rect 422 -223 663 -197
rect 422 -229 664 -223
rect 422 -264 663 -229
rect 422 -268 488 -264
rect 490 -268 660 -264
rect 662 -268 663 -264
rect 422 -282 663 -268
rect 665 -282 706 -171
rect 708 -282 836 -145
rect 460 -283 469 -282
<< nwell >>
rect -1 254 841 299
rect -1 110 841 190
rect -1 1 841 46
rect 2 -2 841 1
rect 417 -34 841 -2
rect 417 -178 841 -98
rect 417 -287 841 -242
<< pwell >>
rect -1 190 841 254
rect -1 46 841 110
rect 417 -98 841 -34
rect 417 -242 841 -178
<< poly >>
rect 13 281 15 286
rect 23 281 25 286
rect 93 288 95 292
rect 33 279 35 283
rect 53 281 55 286
rect 63 281 65 286
rect 13 265 15 268
rect 9 263 15 265
rect 9 261 11 263
rect 13 261 15 263
rect 9 259 15 261
rect 13 246 15 259
rect 23 257 25 268
rect 73 279 75 283
rect 53 265 55 268
rect 49 263 55 265
rect 49 261 51 263
rect 53 261 55 263
rect 33 257 35 261
rect 49 259 55 261
rect 19 255 25 257
rect 19 253 21 255
rect 23 253 25 255
rect 19 251 25 253
rect 29 255 35 257
rect 29 253 31 255
rect 33 253 35 255
rect 29 251 35 253
rect 20 246 22 251
rect 33 246 35 251
rect 53 246 55 259
rect 63 257 65 268
rect 116 285 118 290
rect 123 285 125 290
rect 141 288 143 292
rect 151 288 153 292
rect 161 288 163 292
rect 183 288 185 292
rect 193 288 195 292
rect 203 288 205 292
rect 106 276 108 281
rect 73 257 75 261
rect 59 255 65 257
rect 59 253 61 255
rect 63 253 65 255
rect 59 251 65 253
rect 69 255 75 257
rect 69 253 71 255
rect 73 253 75 255
rect 69 251 75 253
rect 60 246 62 251
rect 73 246 75 251
rect 93 250 95 263
rect 106 260 108 263
rect 221 285 223 290
rect 228 285 230 290
rect 251 288 253 292
rect 272 288 274 292
rect 279 288 281 292
rect 238 276 240 281
rect 360 288 362 292
rect 401 290 403 292
rect 292 278 294 283
rect 320 281 322 286
rect 330 281 332 286
rect 272 264 274 267
rect 238 260 240 263
rect 99 258 108 260
rect 99 256 101 258
rect 103 256 105 258
rect 116 257 118 260
rect 123 257 125 260
rect 141 257 143 260
rect 151 257 153 260
rect 161 257 163 260
rect 183 257 185 260
rect 193 257 195 260
rect 203 257 205 260
rect 221 257 223 260
rect 228 257 230 260
rect 238 258 247 260
rect 99 254 105 256
rect 93 248 99 250
rect 93 246 95 248
rect 97 246 99 248
rect 13 230 15 235
rect 20 230 22 235
rect 33 233 35 237
rect 93 244 99 246
rect 93 241 95 244
rect 103 241 105 254
rect 113 255 119 257
rect 113 253 115 255
rect 117 253 119 255
rect 113 251 119 253
rect 123 255 145 257
rect 123 253 134 255
rect 136 253 141 255
rect 143 253 145 255
rect 123 251 145 253
rect 149 255 155 257
rect 149 253 151 255
rect 153 253 155 255
rect 149 251 155 253
rect 159 255 165 257
rect 159 253 161 255
rect 163 253 165 255
rect 159 251 165 253
rect 181 255 187 257
rect 181 253 183 255
rect 185 253 187 255
rect 181 251 187 253
rect 191 255 197 257
rect 191 253 193 255
rect 195 253 197 255
rect 191 251 197 253
rect 201 255 223 257
rect 201 253 203 255
rect 205 253 210 255
rect 212 253 223 255
rect 201 251 223 253
rect 227 255 233 257
rect 227 253 229 255
rect 231 253 233 255
rect 227 251 233 253
rect 113 248 115 251
rect 123 248 125 251
rect 143 248 145 251
rect 150 248 152 251
rect 53 230 55 235
rect 60 230 62 235
rect 73 233 75 237
rect 93 224 95 228
rect 103 226 105 231
rect 113 229 115 234
rect 123 229 125 234
rect 161 242 163 251
rect 183 242 185 251
rect 194 248 196 251
rect 201 248 203 251
rect 221 248 223 251
rect 231 248 233 251
rect 241 256 243 258
rect 245 256 247 258
rect 241 254 247 256
rect 241 241 243 254
rect 251 250 253 263
rect 268 262 274 264
rect 268 260 270 262
rect 272 260 274 262
rect 268 258 274 260
rect 247 248 253 250
rect 272 248 274 258
rect 279 257 281 267
rect 340 279 342 283
rect 320 265 322 268
rect 316 263 322 265
rect 316 261 318 263
rect 320 261 322 263
rect 292 257 294 260
rect 316 259 322 261
rect 278 255 284 257
rect 278 253 280 255
rect 282 253 284 255
rect 278 251 284 253
rect 288 255 294 257
rect 288 253 290 255
rect 292 253 294 255
rect 288 251 294 253
rect 282 248 284 251
rect 292 248 294 251
rect 247 246 249 248
rect 251 246 253 248
rect 247 244 253 246
rect 251 241 253 244
rect 221 229 223 234
rect 231 229 233 234
rect 143 224 145 228
rect 150 224 152 228
rect 161 224 163 228
rect 183 224 185 228
rect 194 224 196 228
rect 201 224 203 228
rect 241 226 243 231
rect 272 237 274 242
rect 282 237 284 242
rect 320 246 322 259
rect 330 257 332 268
rect 383 285 385 290
rect 390 285 392 290
rect 408 288 410 292
rect 418 288 420 292
rect 428 288 430 292
rect 450 288 452 292
rect 460 288 462 292
rect 470 288 472 292
rect 373 276 375 281
rect 340 257 342 261
rect 326 255 332 257
rect 326 253 328 255
rect 330 253 332 255
rect 326 251 332 253
rect 336 255 342 257
rect 336 253 338 255
rect 340 253 342 255
rect 336 251 342 253
rect 327 246 329 251
rect 340 246 342 251
rect 360 250 362 263
rect 373 260 375 263
rect 488 285 490 290
rect 495 285 497 290
rect 518 288 520 292
rect 539 288 541 292
rect 546 288 548 292
rect 586 290 588 292
rect 505 276 507 281
rect 627 288 629 292
rect 559 278 561 283
rect 587 281 589 286
rect 597 281 599 286
rect 539 264 541 267
rect 505 260 507 263
rect 366 258 375 260
rect 366 256 368 258
rect 370 256 372 258
rect 383 257 385 260
rect 390 257 392 260
rect 408 257 410 260
rect 418 257 420 260
rect 428 257 430 260
rect 450 257 452 260
rect 460 257 462 260
rect 470 257 472 260
rect 488 257 490 260
rect 495 257 497 260
rect 505 258 514 260
rect 366 254 372 256
rect 360 248 366 250
rect 360 246 362 248
rect 364 246 366 248
rect 292 234 294 239
rect 360 244 366 246
rect 360 241 362 244
rect 370 241 372 254
rect 380 255 386 257
rect 380 253 382 255
rect 384 253 386 255
rect 380 251 386 253
rect 390 255 412 257
rect 390 253 401 255
rect 403 253 408 255
rect 410 253 412 255
rect 390 251 412 253
rect 416 255 422 257
rect 416 253 418 255
rect 420 253 422 255
rect 416 251 422 253
rect 426 255 432 257
rect 426 253 428 255
rect 430 253 432 255
rect 426 251 432 253
rect 448 255 454 257
rect 448 253 450 255
rect 452 253 454 255
rect 448 251 454 253
rect 458 255 464 257
rect 458 253 460 255
rect 462 253 464 255
rect 458 251 464 253
rect 468 255 490 257
rect 468 253 470 255
rect 472 253 477 255
rect 479 253 490 255
rect 468 251 490 253
rect 494 255 500 257
rect 494 253 496 255
rect 498 253 500 255
rect 494 251 500 253
rect 380 248 382 251
rect 390 248 392 251
rect 410 248 412 251
rect 417 248 419 251
rect 320 230 322 235
rect 327 230 329 235
rect 251 224 253 228
rect 340 233 342 237
rect 360 224 362 228
rect 370 226 372 231
rect 380 229 382 234
rect 390 229 392 234
rect 428 242 430 251
rect 450 242 452 251
rect 461 248 463 251
rect 468 248 470 251
rect 488 248 490 251
rect 498 248 500 251
rect 508 256 510 258
rect 512 256 514 258
rect 508 254 514 256
rect 508 241 510 254
rect 518 250 520 263
rect 535 262 541 264
rect 535 260 537 262
rect 539 260 541 262
rect 535 258 541 260
rect 514 248 520 250
rect 539 248 541 258
rect 546 257 548 267
rect 607 279 609 283
rect 587 265 589 268
rect 583 263 589 265
rect 583 261 585 263
rect 587 261 589 263
rect 559 257 561 260
rect 583 259 589 261
rect 545 255 551 257
rect 545 253 547 255
rect 549 253 551 255
rect 545 251 551 253
rect 555 255 561 257
rect 555 253 557 255
rect 559 253 561 255
rect 555 251 561 253
rect 549 248 551 251
rect 559 248 561 251
rect 514 246 516 248
rect 518 246 520 248
rect 514 244 520 246
rect 518 241 520 244
rect 488 229 490 234
rect 498 229 500 234
rect 410 224 412 228
rect 417 224 419 228
rect 428 224 430 228
rect 450 224 452 228
rect 461 224 463 228
rect 468 224 470 228
rect 508 226 510 231
rect 539 237 541 242
rect 549 237 551 242
rect 587 246 589 259
rect 597 257 599 268
rect 650 285 652 290
rect 657 285 659 290
rect 675 288 677 292
rect 685 288 687 292
rect 695 288 697 292
rect 717 288 719 292
rect 727 288 729 292
rect 737 288 739 292
rect 778 290 780 292
rect 640 276 642 281
rect 607 257 609 261
rect 593 255 599 257
rect 593 253 595 255
rect 597 253 599 255
rect 593 251 599 253
rect 603 255 609 257
rect 603 253 605 255
rect 607 253 609 255
rect 603 251 609 253
rect 594 246 596 251
rect 607 246 609 251
rect 627 250 629 263
rect 640 260 642 263
rect 755 285 757 290
rect 762 285 764 290
rect 785 288 787 292
rect 806 288 808 292
rect 813 288 815 292
rect 772 276 774 281
rect 826 278 828 283
rect 806 264 808 267
rect 772 260 774 263
rect 633 258 642 260
rect 633 256 635 258
rect 637 256 639 258
rect 650 257 652 260
rect 657 257 659 260
rect 675 257 677 260
rect 685 257 687 260
rect 695 257 697 260
rect 717 257 719 260
rect 727 257 729 260
rect 737 257 739 260
rect 755 257 757 260
rect 762 257 764 260
rect 772 258 781 260
rect 633 254 639 256
rect 627 248 633 250
rect 627 246 629 248
rect 631 246 633 248
rect 559 234 561 239
rect 627 244 633 246
rect 627 241 629 244
rect 637 241 639 254
rect 647 255 653 257
rect 647 253 649 255
rect 651 253 653 255
rect 647 251 653 253
rect 657 255 679 257
rect 657 253 668 255
rect 670 253 675 255
rect 677 253 679 255
rect 657 251 679 253
rect 683 255 689 257
rect 683 253 685 255
rect 687 253 689 255
rect 683 251 689 253
rect 693 255 699 257
rect 693 253 695 255
rect 697 253 699 255
rect 693 251 699 253
rect 715 255 721 257
rect 715 253 717 255
rect 719 253 721 255
rect 715 251 721 253
rect 725 255 731 257
rect 725 253 727 255
rect 729 253 731 255
rect 725 251 731 253
rect 735 255 757 257
rect 735 253 737 255
rect 739 253 744 255
rect 746 253 757 255
rect 735 251 757 253
rect 761 255 767 257
rect 761 253 763 255
rect 765 253 767 255
rect 761 251 767 253
rect 647 248 649 251
rect 657 248 659 251
rect 677 248 679 251
rect 684 248 686 251
rect 587 230 589 235
rect 594 230 596 235
rect 518 224 520 228
rect 607 233 609 237
rect 627 224 629 228
rect 637 226 639 231
rect 647 229 649 234
rect 657 229 659 234
rect 695 242 697 251
rect 717 242 719 251
rect 728 248 730 251
rect 735 248 737 251
rect 755 248 757 251
rect 765 248 767 251
rect 775 256 777 258
rect 779 256 781 258
rect 775 254 781 256
rect 775 241 777 254
rect 785 250 787 263
rect 802 262 808 264
rect 802 260 804 262
rect 806 260 808 262
rect 802 258 808 260
rect 781 248 787 250
rect 806 248 808 258
rect 813 257 815 267
rect 826 257 828 260
rect 812 255 818 257
rect 812 253 814 255
rect 816 253 818 255
rect 812 251 818 253
rect 822 255 828 257
rect 822 253 824 255
rect 826 253 828 255
rect 822 251 828 253
rect 816 248 818 251
rect 826 248 828 251
rect 781 246 783 248
rect 785 246 787 248
rect 781 244 787 246
rect 785 241 787 244
rect 755 229 757 234
rect 765 229 767 234
rect 677 224 679 228
rect 684 224 686 228
rect 695 224 697 228
rect 717 224 719 228
rect 728 224 730 228
rect 735 224 737 228
rect 775 226 777 231
rect 806 237 808 242
rect 816 237 818 242
rect 826 234 828 239
rect 785 224 787 228
rect 13 209 15 214
rect 20 209 22 214
rect 33 207 35 211
rect 53 209 55 214
rect 60 209 62 214
rect 93 216 95 220
rect 73 207 75 211
rect 103 213 105 218
rect 143 216 145 220
rect 150 216 152 220
rect 161 216 163 220
rect 183 216 185 220
rect 194 216 196 220
rect 201 216 203 220
rect 113 210 115 215
rect 123 210 125 215
rect 93 200 95 203
rect 93 198 99 200
rect 13 185 15 198
rect 20 193 22 198
rect 33 193 35 198
rect 19 191 25 193
rect 19 189 21 191
rect 23 189 25 191
rect 19 187 25 189
rect 29 191 35 193
rect 29 189 31 191
rect 33 189 35 191
rect 29 187 35 189
rect 9 183 15 185
rect 9 181 11 183
rect 13 181 15 183
rect 9 179 15 181
rect 13 176 15 179
rect 23 176 25 187
rect 33 183 35 187
rect 53 185 55 198
rect 60 193 62 198
rect 73 193 75 198
rect 59 191 65 193
rect 59 189 61 191
rect 63 189 65 191
rect 59 187 65 189
rect 69 191 75 193
rect 69 189 71 191
rect 73 189 75 191
rect 69 187 75 189
rect 49 183 55 185
rect 49 181 51 183
rect 53 181 55 183
rect 49 179 55 181
rect 53 176 55 179
rect 63 176 65 187
rect 73 183 75 187
rect 93 196 95 198
rect 97 196 99 198
rect 93 194 99 196
rect 13 158 15 163
rect 23 158 25 163
rect 33 161 35 165
rect 93 181 95 194
rect 103 190 105 203
rect 99 188 105 190
rect 99 186 101 188
rect 103 186 105 188
rect 113 193 115 196
rect 123 193 125 196
rect 143 193 145 196
rect 150 193 152 196
rect 161 193 163 202
rect 183 193 185 202
rect 221 210 223 215
rect 231 210 233 215
rect 241 213 243 218
rect 251 216 253 220
rect 194 193 196 196
rect 201 193 203 196
rect 221 193 223 196
rect 231 193 233 196
rect 113 191 119 193
rect 113 189 115 191
rect 117 189 119 191
rect 113 187 119 189
rect 123 191 145 193
rect 123 189 134 191
rect 136 189 141 191
rect 143 189 145 191
rect 123 187 145 189
rect 149 191 155 193
rect 149 189 151 191
rect 153 189 155 191
rect 149 187 155 189
rect 159 191 165 193
rect 159 189 161 191
rect 163 189 165 191
rect 159 187 165 189
rect 181 191 187 193
rect 181 189 183 191
rect 185 189 187 191
rect 181 187 187 189
rect 191 191 197 193
rect 191 189 193 191
rect 195 189 197 191
rect 191 187 197 189
rect 201 191 223 193
rect 201 189 203 191
rect 205 189 210 191
rect 212 189 223 191
rect 201 187 223 189
rect 227 191 233 193
rect 227 189 229 191
rect 231 189 233 191
rect 227 187 233 189
rect 241 190 243 203
rect 251 200 253 203
rect 247 198 253 200
rect 247 196 249 198
rect 251 196 253 198
rect 272 202 274 207
rect 282 202 284 207
rect 292 205 294 210
rect 320 209 322 214
rect 327 209 329 214
rect 360 216 362 220
rect 340 207 342 211
rect 370 213 372 218
rect 410 216 412 220
rect 417 216 419 220
rect 428 216 430 220
rect 450 216 452 220
rect 461 216 463 220
rect 468 216 470 220
rect 380 210 382 215
rect 390 210 392 215
rect 360 200 362 203
rect 360 198 366 200
rect 247 194 253 196
rect 241 188 247 190
rect 99 184 108 186
rect 116 184 118 187
rect 123 184 125 187
rect 141 184 143 187
rect 151 184 153 187
rect 161 184 163 187
rect 183 184 185 187
rect 193 184 195 187
rect 203 184 205 187
rect 221 184 223 187
rect 228 184 230 187
rect 241 186 243 188
rect 245 186 247 188
rect 238 184 247 186
rect 106 181 108 184
rect 53 158 55 163
rect 63 158 65 163
rect 73 161 75 165
rect 106 163 108 168
rect 93 152 95 156
rect 116 154 118 159
rect 123 154 125 159
rect 238 181 240 184
rect 251 181 253 194
rect 272 186 274 196
rect 282 193 284 196
rect 292 193 294 196
rect 278 191 284 193
rect 278 189 280 191
rect 282 189 284 191
rect 278 187 284 189
rect 288 191 294 193
rect 288 189 290 191
rect 292 189 294 191
rect 288 187 294 189
rect 268 184 274 186
rect 268 182 270 184
rect 272 182 274 184
rect 238 163 240 168
rect 141 152 143 156
rect 151 152 153 156
rect 161 152 163 156
rect 183 152 185 156
rect 193 152 195 156
rect 203 152 205 156
rect 221 154 223 159
rect 228 154 230 159
rect 268 180 274 182
rect 272 177 274 180
rect 279 177 281 187
rect 292 184 294 187
rect 320 185 322 198
rect 327 193 329 198
rect 340 193 342 198
rect 326 191 332 193
rect 326 189 328 191
rect 330 189 332 191
rect 326 187 332 189
rect 336 191 342 193
rect 336 189 338 191
rect 340 189 342 191
rect 336 187 342 189
rect 316 183 322 185
rect 316 181 318 183
rect 320 181 322 183
rect 316 179 322 181
rect 320 176 322 179
rect 330 176 332 187
rect 340 183 342 187
rect 360 196 362 198
rect 364 196 366 198
rect 360 194 366 196
rect 292 161 294 166
rect 360 181 362 194
rect 370 190 372 203
rect 366 188 372 190
rect 366 186 368 188
rect 370 186 372 188
rect 380 193 382 196
rect 390 193 392 196
rect 410 193 412 196
rect 417 193 419 196
rect 428 193 430 202
rect 450 193 452 202
rect 488 210 490 215
rect 498 210 500 215
rect 508 213 510 218
rect 518 216 520 220
rect 461 193 463 196
rect 468 193 470 196
rect 488 193 490 196
rect 498 193 500 196
rect 380 191 386 193
rect 380 189 382 191
rect 384 189 386 191
rect 380 187 386 189
rect 390 191 412 193
rect 390 189 401 191
rect 403 189 408 191
rect 410 189 412 191
rect 390 187 412 189
rect 416 191 422 193
rect 416 189 418 191
rect 420 189 422 191
rect 416 187 422 189
rect 426 191 432 193
rect 426 189 428 191
rect 430 189 432 191
rect 426 187 432 189
rect 448 191 454 193
rect 448 189 450 191
rect 452 189 454 191
rect 448 187 454 189
rect 458 191 464 193
rect 458 189 460 191
rect 462 189 464 191
rect 458 187 464 189
rect 468 191 490 193
rect 468 189 470 191
rect 472 189 477 191
rect 479 189 490 191
rect 468 187 490 189
rect 494 191 500 193
rect 494 189 496 191
rect 498 189 500 191
rect 494 187 500 189
rect 508 190 510 203
rect 518 200 520 203
rect 514 198 520 200
rect 514 196 516 198
rect 518 196 520 198
rect 539 202 541 207
rect 549 202 551 207
rect 559 205 561 210
rect 587 209 589 214
rect 594 209 596 214
rect 627 216 629 220
rect 607 207 609 211
rect 637 213 639 218
rect 677 216 679 220
rect 684 216 686 220
rect 695 216 697 220
rect 717 216 719 220
rect 728 216 730 220
rect 735 216 737 220
rect 647 210 649 215
rect 657 210 659 215
rect 627 200 629 203
rect 627 198 633 200
rect 514 194 520 196
rect 508 188 514 190
rect 366 184 375 186
rect 383 184 385 187
rect 390 184 392 187
rect 408 184 410 187
rect 418 184 420 187
rect 428 184 430 187
rect 450 184 452 187
rect 460 184 462 187
rect 470 184 472 187
rect 488 184 490 187
rect 495 184 497 187
rect 508 186 510 188
rect 512 186 514 188
rect 505 184 514 186
rect 373 181 375 184
rect 320 158 322 163
rect 330 158 332 163
rect 340 161 342 165
rect 251 152 253 156
rect 272 152 274 156
rect 279 152 281 156
rect 373 163 375 168
rect 360 152 362 156
rect 383 154 385 159
rect 390 154 392 159
rect 505 181 507 184
rect 518 181 520 194
rect 539 186 541 196
rect 549 193 551 196
rect 559 193 561 196
rect 545 191 551 193
rect 545 189 547 191
rect 549 189 551 191
rect 545 187 551 189
rect 555 191 561 193
rect 555 189 557 191
rect 559 189 561 191
rect 555 187 561 189
rect 535 184 541 186
rect 535 182 537 184
rect 539 182 541 184
rect 505 163 507 168
rect 408 152 410 156
rect 418 152 420 156
rect 428 152 430 156
rect 450 152 452 156
rect 460 152 462 156
rect 470 152 472 156
rect 488 154 490 159
rect 495 154 497 159
rect 535 180 541 182
rect 539 177 541 180
rect 546 177 548 187
rect 559 184 561 187
rect 587 185 589 198
rect 594 193 596 198
rect 607 193 609 198
rect 593 191 599 193
rect 593 189 595 191
rect 597 189 599 191
rect 593 187 599 189
rect 603 191 609 193
rect 603 189 605 191
rect 607 189 609 191
rect 603 187 609 189
rect 583 183 589 185
rect 583 181 585 183
rect 587 181 589 183
rect 583 179 589 181
rect 587 176 589 179
rect 597 176 599 187
rect 607 183 609 187
rect 627 196 629 198
rect 631 196 633 198
rect 627 194 633 196
rect 559 161 561 166
rect 627 181 629 194
rect 637 190 639 203
rect 633 188 639 190
rect 633 186 635 188
rect 637 186 639 188
rect 647 193 649 196
rect 657 193 659 196
rect 677 193 679 196
rect 684 193 686 196
rect 695 193 697 202
rect 717 193 719 202
rect 755 210 757 215
rect 765 210 767 215
rect 775 213 777 218
rect 785 216 787 220
rect 728 193 730 196
rect 735 193 737 196
rect 755 193 757 196
rect 765 193 767 196
rect 647 191 653 193
rect 647 189 649 191
rect 651 189 653 191
rect 647 187 653 189
rect 657 191 679 193
rect 657 189 668 191
rect 670 189 675 191
rect 677 189 679 191
rect 657 187 679 189
rect 683 191 689 193
rect 683 189 685 191
rect 687 189 689 191
rect 683 187 689 189
rect 693 191 699 193
rect 693 189 695 191
rect 697 189 699 191
rect 693 187 699 189
rect 715 191 721 193
rect 715 189 717 191
rect 719 189 721 191
rect 715 187 721 189
rect 725 191 731 193
rect 725 189 727 191
rect 729 189 731 191
rect 725 187 731 189
rect 735 191 757 193
rect 735 189 737 191
rect 739 189 744 191
rect 746 189 757 191
rect 735 187 757 189
rect 761 191 767 193
rect 761 189 763 191
rect 765 189 767 191
rect 761 187 767 189
rect 775 190 777 203
rect 785 200 787 203
rect 781 198 787 200
rect 781 196 783 198
rect 785 196 787 198
rect 806 202 808 207
rect 816 202 818 207
rect 826 205 828 210
rect 781 194 787 196
rect 775 188 781 190
rect 633 184 642 186
rect 650 184 652 187
rect 657 184 659 187
rect 675 184 677 187
rect 685 184 687 187
rect 695 184 697 187
rect 717 184 719 187
rect 727 184 729 187
rect 737 184 739 187
rect 755 184 757 187
rect 762 184 764 187
rect 775 186 777 188
rect 779 186 781 188
rect 772 184 781 186
rect 640 181 642 184
rect 587 158 589 163
rect 597 158 599 163
rect 607 161 609 165
rect 518 152 520 156
rect 539 152 541 156
rect 546 152 548 156
rect 640 163 642 168
rect 627 152 629 156
rect 650 154 652 159
rect 657 154 659 159
rect 772 181 774 184
rect 785 181 787 194
rect 806 186 808 196
rect 816 193 818 196
rect 826 193 828 196
rect 812 191 818 193
rect 812 189 814 191
rect 816 189 818 191
rect 812 187 818 189
rect 822 191 828 193
rect 822 189 824 191
rect 826 189 828 191
rect 822 187 828 189
rect 802 184 808 186
rect 802 182 804 184
rect 806 182 808 184
rect 772 163 774 168
rect 675 152 677 156
rect 685 152 687 156
rect 695 152 697 156
rect 717 152 719 156
rect 727 152 729 156
rect 737 152 739 156
rect 755 154 757 159
rect 762 154 764 159
rect 802 180 808 182
rect 806 177 808 180
rect 813 177 815 187
rect 826 184 828 187
rect 826 161 828 166
rect 785 152 787 156
rect 806 152 808 156
rect 813 152 815 156
rect 832 149 834 151
rect 13 137 15 142
rect 23 137 25 142
rect 93 144 95 148
rect 33 135 35 139
rect 53 137 55 142
rect 63 137 65 142
rect 13 121 15 124
rect 9 119 15 121
rect 9 117 11 119
rect 13 117 15 119
rect 9 115 15 117
rect 13 102 15 115
rect 23 113 25 124
rect 73 135 75 139
rect 53 121 55 124
rect 49 119 55 121
rect 49 117 51 119
rect 53 117 55 119
rect 33 113 35 117
rect 49 115 55 117
rect 19 111 25 113
rect 19 109 21 111
rect 23 109 25 111
rect 19 107 25 109
rect 29 111 35 113
rect 29 109 31 111
rect 33 109 35 111
rect 29 107 35 109
rect 20 102 22 107
rect 33 102 35 107
rect 53 102 55 115
rect 63 113 65 124
rect 116 141 118 146
rect 123 141 125 146
rect 141 144 143 148
rect 151 144 153 148
rect 161 144 163 148
rect 183 144 185 148
rect 193 144 195 148
rect 203 144 205 148
rect 106 132 108 137
rect 73 113 75 117
rect 59 111 65 113
rect 59 109 61 111
rect 63 109 65 111
rect 59 107 65 109
rect 69 111 75 113
rect 69 109 71 111
rect 73 109 75 111
rect 69 107 75 109
rect 60 102 62 107
rect 73 102 75 107
rect 93 106 95 119
rect 106 116 108 119
rect 221 141 223 146
rect 228 141 230 146
rect 251 144 253 148
rect 272 144 274 148
rect 279 144 281 148
rect 238 132 240 137
rect 360 144 362 148
rect 292 134 294 139
rect 320 137 322 142
rect 330 137 332 142
rect 272 120 274 123
rect 238 116 240 119
rect 99 114 108 116
rect 99 112 101 114
rect 103 112 105 114
rect 116 113 118 116
rect 123 113 125 116
rect 141 113 143 116
rect 151 113 153 116
rect 161 113 163 116
rect 183 113 185 116
rect 193 113 195 116
rect 203 113 205 116
rect 221 113 223 116
rect 228 113 230 116
rect 238 114 247 116
rect 99 110 105 112
rect 93 104 99 106
rect 93 102 95 104
rect 97 102 99 104
rect 13 86 15 91
rect 20 86 22 91
rect 33 89 35 93
rect 93 100 99 102
rect 93 97 95 100
rect 103 97 105 110
rect 113 111 119 113
rect 113 109 115 111
rect 117 109 119 111
rect 113 107 119 109
rect 123 111 145 113
rect 123 109 134 111
rect 136 109 141 111
rect 143 109 145 111
rect 123 107 145 109
rect 149 111 155 113
rect 149 109 151 111
rect 153 109 155 111
rect 149 107 155 109
rect 159 111 165 113
rect 159 109 161 111
rect 163 109 165 111
rect 159 107 165 109
rect 181 111 187 113
rect 181 109 183 111
rect 185 109 187 111
rect 181 107 187 109
rect 191 111 197 113
rect 191 109 193 111
rect 195 109 197 111
rect 191 107 197 109
rect 201 111 223 113
rect 201 109 203 111
rect 205 109 210 111
rect 212 109 223 111
rect 201 107 223 109
rect 227 111 233 113
rect 227 109 229 111
rect 231 109 233 111
rect 227 107 233 109
rect 113 104 115 107
rect 123 104 125 107
rect 143 104 145 107
rect 150 104 152 107
rect 53 86 55 91
rect 60 86 62 91
rect 73 89 75 93
rect 93 80 95 84
rect 103 82 105 87
rect 113 85 115 90
rect 123 85 125 90
rect 161 98 163 107
rect 183 98 185 107
rect 194 104 196 107
rect 201 104 203 107
rect 221 104 223 107
rect 231 104 233 107
rect 241 112 243 114
rect 245 112 247 114
rect 241 110 247 112
rect 241 97 243 110
rect 251 106 253 119
rect 268 118 274 120
rect 268 116 270 118
rect 272 116 274 118
rect 268 114 274 116
rect 247 104 253 106
rect 272 104 274 114
rect 279 113 281 123
rect 340 135 342 139
rect 320 121 322 124
rect 316 119 322 121
rect 316 117 318 119
rect 320 117 322 119
rect 292 113 294 116
rect 316 115 322 117
rect 278 111 284 113
rect 278 109 280 111
rect 282 109 284 111
rect 278 107 284 109
rect 288 111 294 113
rect 288 109 290 111
rect 292 109 294 111
rect 288 107 294 109
rect 282 104 284 107
rect 292 104 294 107
rect 247 102 249 104
rect 251 102 253 104
rect 247 100 253 102
rect 251 97 253 100
rect 221 85 223 90
rect 231 85 233 90
rect 143 80 145 84
rect 150 80 152 84
rect 161 80 163 84
rect 183 80 185 84
rect 194 80 196 84
rect 201 80 203 84
rect 241 82 243 87
rect 272 93 274 98
rect 282 93 284 98
rect 320 102 322 115
rect 330 113 332 124
rect 383 141 385 146
rect 390 141 392 146
rect 408 144 410 148
rect 418 144 420 148
rect 428 144 430 148
rect 450 144 452 148
rect 460 144 462 148
rect 470 144 472 148
rect 373 132 375 137
rect 340 113 342 117
rect 326 111 332 113
rect 326 109 328 111
rect 330 109 332 111
rect 326 107 332 109
rect 336 111 342 113
rect 336 109 338 111
rect 340 109 342 111
rect 336 107 342 109
rect 327 102 329 107
rect 340 102 342 107
rect 360 106 362 119
rect 373 116 375 119
rect 488 141 490 146
rect 495 141 497 146
rect 518 144 520 148
rect 539 144 541 148
rect 546 144 548 148
rect 505 132 507 137
rect 627 144 629 148
rect 559 134 561 139
rect 587 137 589 142
rect 597 137 599 142
rect 539 120 541 123
rect 505 116 507 119
rect 366 114 375 116
rect 366 112 368 114
rect 370 112 372 114
rect 383 113 385 116
rect 390 113 392 116
rect 408 113 410 116
rect 418 113 420 116
rect 428 113 430 116
rect 450 113 452 116
rect 460 113 462 116
rect 470 113 472 116
rect 488 113 490 116
rect 495 113 497 116
rect 505 114 514 116
rect 366 110 372 112
rect 360 104 366 106
rect 360 102 362 104
rect 364 102 366 104
rect 292 90 294 95
rect 360 100 366 102
rect 360 97 362 100
rect 370 97 372 110
rect 380 111 386 113
rect 380 109 382 111
rect 384 109 386 111
rect 380 107 386 109
rect 390 111 412 113
rect 390 109 401 111
rect 403 109 408 111
rect 410 109 412 111
rect 390 107 412 109
rect 416 111 422 113
rect 416 109 418 111
rect 420 109 422 111
rect 416 107 422 109
rect 426 111 432 113
rect 426 109 428 111
rect 430 109 432 111
rect 426 107 432 109
rect 448 111 454 113
rect 448 109 450 111
rect 452 109 454 111
rect 448 107 454 109
rect 458 111 464 113
rect 458 109 460 111
rect 462 109 464 111
rect 458 107 464 109
rect 468 111 490 113
rect 468 109 470 111
rect 472 109 477 111
rect 479 109 490 111
rect 468 107 490 109
rect 494 111 500 113
rect 494 109 496 111
rect 498 109 500 111
rect 494 107 500 109
rect 380 104 382 107
rect 390 104 392 107
rect 410 104 412 107
rect 417 104 419 107
rect 320 86 322 91
rect 327 86 329 91
rect 251 80 253 84
rect 340 89 342 93
rect 360 80 362 84
rect 370 82 372 87
rect 380 85 382 90
rect 390 85 392 90
rect 428 98 430 107
rect 450 98 452 107
rect 461 104 463 107
rect 468 104 470 107
rect 488 104 490 107
rect 498 104 500 107
rect 508 112 510 114
rect 512 112 514 114
rect 508 110 514 112
rect 508 97 510 110
rect 518 106 520 119
rect 535 118 541 120
rect 535 116 537 118
rect 539 116 541 118
rect 535 114 541 116
rect 514 104 520 106
rect 539 104 541 114
rect 546 113 548 123
rect 607 135 609 139
rect 587 121 589 124
rect 583 119 589 121
rect 583 117 585 119
rect 587 117 589 119
rect 559 113 561 116
rect 583 115 589 117
rect 545 111 551 113
rect 545 109 547 111
rect 549 109 551 111
rect 545 107 551 109
rect 555 111 561 113
rect 555 109 557 111
rect 559 109 561 111
rect 555 107 561 109
rect 549 104 551 107
rect 559 104 561 107
rect 514 102 516 104
rect 518 102 520 104
rect 514 100 520 102
rect 518 97 520 100
rect 488 85 490 90
rect 498 85 500 90
rect 410 80 412 84
rect 417 80 419 84
rect 428 80 430 84
rect 450 80 452 84
rect 461 80 463 84
rect 468 80 470 84
rect 508 82 510 87
rect 539 93 541 98
rect 549 93 551 98
rect 587 102 589 115
rect 597 113 599 124
rect 650 141 652 146
rect 657 141 659 146
rect 675 144 677 148
rect 685 144 687 148
rect 695 144 697 148
rect 717 144 719 148
rect 727 144 729 148
rect 737 144 739 148
rect 640 132 642 137
rect 607 113 609 117
rect 593 111 599 113
rect 593 109 595 111
rect 597 109 599 111
rect 593 107 599 109
rect 603 111 609 113
rect 603 109 605 111
rect 607 109 609 111
rect 603 107 609 109
rect 594 102 596 107
rect 607 102 609 107
rect 627 106 629 119
rect 640 116 642 119
rect 755 141 757 146
rect 762 141 764 146
rect 785 144 787 148
rect 806 144 808 148
rect 813 144 815 148
rect 772 132 774 137
rect 826 134 828 139
rect 806 120 808 123
rect 772 116 774 119
rect 633 114 642 116
rect 633 112 635 114
rect 637 112 639 114
rect 650 113 652 116
rect 657 113 659 116
rect 675 113 677 116
rect 685 113 687 116
rect 695 113 697 116
rect 717 113 719 116
rect 727 113 729 116
rect 737 113 739 116
rect 755 113 757 116
rect 762 113 764 116
rect 772 114 781 116
rect 633 110 639 112
rect 627 104 633 106
rect 627 102 629 104
rect 631 102 633 104
rect 559 90 561 95
rect 627 100 633 102
rect 627 97 629 100
rect 637 97 639 110
rect 647 111 653 113
rect 647 109 649 111
rect 651 109 653 111
rect 647 107 653 109
rect 657 111 679 113
rect 657 109 668 111
rect 670 109 675 111
rect 677 109 679 111
rect 657 107 679 109
rect 683 111 689 113
rect 683 109 685 111
rect 687 109 689 111
rect 683 107 689 109
rect 693 111 699 113
rect 693 109 695 111
rect 697 109 699 111
rect 693 107 699 109
rect 715 111 721 113
rect 715 109 717 111
rect 719 109 721 111
rect 715 107 721 109
rect 725 111 731 113
rect 725 109 727 111
rect 729 109 731 111
rect 725 107 731 109
rect 735 111 757 113
rect 735 109 737 111
rect 739 109 744 111
rect 746 109 757 111
rect 735 107 757 109
rect 761 111 767 113
rect 761 109 763 111
rect 765 109 767 111
rect 761 107 767 109
rect 647 104 649 107
rect 657 104 659 107
rect 677 104 679 107
rect 684 104 686 107
rect 587 86 589 91
rect 594 86 596 91
rect 518 80 520 84
rect 607 89 609 93
rect 627 80 629 84
rect 637 82 639 87
rect 647 85 649 90
rect 657 85 659 90
rect 695 98 697 107
rect 717 98 719 107
rect 728 104 730 107
rect 735 104 737 107
rect 755 104 757 107
rect 765 104 767 107
rect 775 112 777 114
rect 779 112 781 114
rect 775 110 781 112
rect 775 97 777 110
rect 785 106 787 119
rect 802 118 808 120
rect 802 116 804 118
rect 806 116 808 118
rect 802 114 808 116
rect 781 104 787 106
rect 806 104 808 114
rect 813 113 815 123
rect 826 113 828 116
rect 812 111 818 113
rect 812 109 814 111
rect 816 109 818 111
rect 812 107 818 109
rect 822 111 828 113
rect 822 109 824 111
rect 826 109 828 111
rect 822 107 828 109
rect 816 104 818 107
rect 826 104 828 107
rect 781 102 783 104
rect 785 102 787 104
rect 781 100 787 102
rect 785 97 787 100
rect 755 85 757 90
rect 765 85 767 90
rect 677 80 679 84
rect 684 80 686 84
rect 695 80 697 84
rect 717 80 719 84
rect 728 80 730 84
rect 735 80 737 84
rect 775 82 777 87
rect 806 93 808 98
rect 816 93 818 98
rect 826 90 828 95
rect 785 80 787 84
rect 13 65 15 70
rect 20 65 22 70
rect 33 63 35 67
rect 53 65 55 70
rect 60 65 62 70
rect 93 72 95 76
rect 73 63 75 67
rect 103 69 105 74
rect 143 72 145 76
rect 150 72 152 76
rect 161 72 163 76
rect 183 72 185 76
rect 194 72 196 76
rect 201 72 203 76
rect 113 66 115 71
rect 123 66 125 71
rect 93 56 95 59
rect 93 54 99 56
rect 13 41 15 54
rect 20 49 22 54
rect 33 49 35 54
rect 19 47 25 49
rect 19 45 21 47
rect 23 45 25 47
rect 19 43 25 45
rect 29 47 35 49
rect 29 45 31 47
rect 33 45 35 47
rect 29 43 35 45
rect 9 39 15 41
rect 9 37 11 39
rect 13 37 15 39
rect 9 35 15 37
rect 13 32 15 35
rect 23 32 25 43
rect 33 39 35 43
rect 53 41 55 54
rect 60 49 62 54
rect 73 49 75 54
rect 59 47 65 49
rect 59 45 61 47
rect 63 45 65 47
rect 59 43 65 45
rect 69 47 75 49
rect 69 45 71 47
rect 73 45 75 47
rect 69 43 75 45
rect 49 39 55 41
rect 49 37 51 39
rect 53 37 55 39
rect 49 35 55 37
rect 53 32 55 35
rect 63 32 65 43
rect 73 39 75 43
rect 93 52 95 54
rect 97 52 99 54
rect 93 50 99 52
rect 13 14 15 19
rect 23 14 25 19
rect 33 17 35 21
rect 93 37 95 50
rect 103 46 105 59
rect 99 44 105 46
rect 99 42 101 44
rect 103 42 105 44
rect 113 49 115 52
rect 123 49 125 52
rect 143 49 145 52
rect 150 49 152 52
rect 161 49 163 58
rect 183 49 185 58
rect 221 66 223 71
rect 231 66 233 71
rect 241 69 243 74
rect 251 72 253 76
rect 194 49 196 52
rect 201 49 203 52
rect 221 49 223 52
rect 231 49 233 52
rect 113 47 119 49
rect 113 45 115 47
rect 117 45 119 47
rect 113 43 119 45
rect 123 47 145 49
rect 123 45 134 47
rect 136 45 141 47
rect 143 45 145 47
rect 123 43 145 45
rect 149 47 155 49
rect 149 45 151 47
rect 153 45 155 47
rect 149 43 155 45
rect 159 47 165 49
rect 159 45 161 47
rect 163 45 165 47
rect 159 43 165 45
rect 181 47 187 49
rect 181 45 183 47
rect 185 45 187 47
rect 181 43 187 45
rect 191 47 197 49
rect 191 45 193 47
rect 195 45 197 47
rect 191 43 197 45
rect 201 47 223 49
rect 201 45 203 47
rect 205 45 210 47
rect 212 45 223 47
rect 201 43 223 45
rect 227 47 233 49
rect 227 45 229 47
rect 231 45 233 47
rect 227 43 233 45
rect 241 46 243 59
rect 251 56 253 59
rect 247 54 253 56
rect 247 52 249 54
rect 251 52 253 54
rect 272 58 274 63
rect 282 58 284 63
rect 292 61 294 66
rect 320 65 322 70
rect 327 65 329 70
rect 360 72 362 76
rect 340 63 342 67
rect 370 69 372 74
rect 410 72 412 76
rect 417 72 419 76
rect 428 72 430 76
rect 450 72 452 76
rect 461 72 463 76
rect 468 72 470 76
rect 380 66 382 71
rect 390 66 392 71
rect 360 56 362 59
rect 360 54 366 56
rect 247 50 253 52
rect 241 44 247 46
rect 99 40 108 42
rect 116 40 118 43
rect 123 40 125 43
rect 141 40 143 43
rect 151 40 153 43
rect 161 40 163 43
rect 183 40 185 43
rect 193 40 195 43
rect 203 40 205 43
rect 221 40 223 43
rect 228 40 230 43
rect 241 42 243 44
rect 245 42 247 44
rect 238 40 247 42
rect 106 37 108 40
rect 53 14 55 19
rect 63 14 65 19
rect 73 17 75 21
rect 106 19 108 24
rect 93 8 95 12
rect 116 10 118 15
rect 123 10 125 15
rect 238 37 240 40
rect 251 37 253 50
rect 272 42 274 52
rect 282 49 284 52
rect 292 49 294 52
rect 278 47 284 49
rect 278 45 280 47
rect 282 45 284 47
rect 278 43 284 45
rect 288 47 294 49
rect 288 45 290 47
rect 292 45 294 47
rect 288 43 294 45
rect 268 40 274 42
rect 268 38 270 40
rect 272 38 274 40
rect 238 19 240 24
rect 141 8 143 12
rect 151 8 153 12
rect 161 8 163 12
rect 183 8 185 12
rect 193 8 195 12
rect 203 8 205 12
rect 221 10 223 15
rect 228 10 230 15
rect 268 36 274 38
rect 272 33 274 36
rect 279 33 281 43
rect 292 40 294 43
rect 320 41 322 54
rect 327 49 329 54
rect 340 49 342 54
rect 326 47 332 49
rect 326 45 328 47
rect 330 45 332 47
rect 326 43 332 45
rect 336 47 342 49
rect 336 45 338 47
rect 340 45 342 47
rect 336 43 342 45
rect 316 39 322 41
rect 316 37 318 39
rect 320 37 322 39
rect 316 35 322 37
rect 320 32 322 35
rect 330 32 332 43
rect 340 39 342 43
rect 360 52 362 54
rect 364 52 366 54
rect 360 50 366 52
rect 292 17 294 22
rect 360 37 362 50
rect 370 46 372 59
rect 366 44 372 46
rect 366 42 368 44
rect 370 42 372 44
rect 380 49 382 52
rect 390 49 392 52
rect 410 49 412 52
rect 417 49 419 52
rect 428 49 430 58
rect 450 49 452 58
rect 488 66 490 71
rect 498 66 500 71
rect 508 69 510 74
rect 518 72 520 76
rect 461 49 463 52
rect 468 49 470 52
rect 488 49 490 52
rect 498 49 500 52
rect 380 47 386 49
rect 380 45 382 47
rect 384 45 386 47
rect 380 43 386 45
rect 390 47 412 49
rect 390 45 401 47
rect 403 45 408 47
rect 410 45 412 47
rect 390 43 412 45
rect 416 47 422 49
rect 416 45 418 47
rect 420 45 422 47
rect 416 43 422 45
rect 426 47 432 49
rect 426 45 428 47
rect 430 45 432 47
rect 426 43 432 45
rect 448 47 454 49
rect 448 45 450 47
rect 452 45 454 47
rect 448 43 454 45
rect 458 47 464 49
rect 458 45 460 47
rect 462 45 464 47
rect 458 43 464 45
rect 468 47 490 49
rect 468 45 470 47
rect 472 45 477 47
rect 479 45 490 47
rect 468 43 490 45
rect 494 47 500 49
rect 494 45 496 47
rect 498 45 500 47
rect 494 43 500 45
rect 508 46 510 59
rect 518 56 520 59
rect 514 54 520 56
rect 514 52 516 54
rect 518 52 520 54
rect 539 58 541 63
rect 549 58 551 63
rect 559 61 561 66
rect 587 65 589 70
rect 594 65 596 70
rect 627 72 629 76
rect 607 63 609 67
rect 637 69 639 74
rect 677 72 679 76
rect 684 72 686 76
rect 695 72 697 76
rect 717 72 719 76
rect 728 72 730 76
rect 735 72 737 76
rect 647 66 649 71
rect 657 66 659 71
rect 627 56 629 59
rect 627 54 633 56
rect 514 50 520 52
rect 508 44 514 46
rect 366 40 375 42
rect 383 40 385 43
rect 390 40 392 43
rect 408 40 410 43
rect 418 40 420 43
rect 428 40 430 43
rect 450 40 452 43
rect 460 40 462 43
rect 470 40 472 43
rect 488 40 490 43
rect 495 40 497 43
rect 508 42 510 44
rect 512 42 514 44
rect 505 40 514 42
rect 373 37 375 40
rect 320 14 322 19
rect 330 14 332 19
rect 340 17 342 21
rect 251 8 253 12
rect 272 8 274 12
rect 279 8 281 12
rect 373 19 375 24
rect 360 8 362 12
rect 383 10 385 15
rect 390 10 392 15
rect 505 37 507 40
rect 518 37 520 50
rect 539 42 541 52
rect 549 49 551 52
rect 559 49 561 52
rect 545 47 551 49
rect 545 45 547 47
rect 549 45 551 47
rect 545 43 551 45
rect 555 47 561 49
rect 555 45 557 47
rect 559 45 561 47
rect 555 43 561 45
rect 535 40 541 42
rect 535 38 537 40
rect 539 38 541 40
rect 505 19 507 24
rect 408 8 410 12
rect 418 8 420 12
rect 428 8 430 12
rect 450 8 452 12
rect 460 8 462 12
rect 470 8 472 12
rect 488 10 490 15
rect 495 10 497 15
rect 535 36 541 38
rect 539 33 541 36
rect 546 33 548 43
rect 559 40 561 43
rect 587 41 589 54
rect 594 49 596 54
rect 607 49 609 54
rect 593 47 599 49
rect 593 45 595 47
rect 597 45 599 47
rect 593 43 599 45
rect 603 47 609 49
rect 603 45 605 47
rect 607 45 609 47
rect 603 43 609 45
rect 583 39 589 41
rect 583 37 585 39
rect 587 37 589 39
rect 583 35 589 37
rect 587 32 589 35
rect 597 32 599 43
rect 607 39 609 43
rect 627 52 629 54
rect 631 52 633 54
rect 627 50 633 52
rect 559 17 561 22
rect 627 37 629 50
rect 637 46 639 59
rect 633 44 639 46
rect 633 42 635 44
rect 637 42 639 44
rect 647 49 649 52
rect 657 49 659 52
rect 677 49 679 52
rect 684 49 686 52
rect 695 49 697 58
rect 717 49 719 58
rect 755 66 757 71
rect 765 66 767 71
rect 775 69 777 74
rect 785 72 787 76
rect 728 49 730 52
rect 735 49 737 52
rect 755 49 757 52
rect 765 49 767 52
rect 647 47 653 49
rect 647 45 649 47
rect 651 45 653 47
rect 647 43 653 45
rect 657 47 679 49
rect 657 45 668 47
rect 670 45 675 47
rect 677 45 679 47
rect 657 43 679 45
rect 683 47 689 49
rect 683 45 685 47
rect 687 45 689 47
rect 683 43 689 45
rect 693 47 699 49
rect 693 45 695 47
rect 697 45 699 47
rect 693 43 699 45
rect 715 47 721 49
rect 715 45 717 47
rect 719 45 721 47
rect 715 43 721 45
rect 725 47 731 49
rect 725 45 727 47
rect 729 45 731 47
rect 725 43 731 45
rect 735 47 757 49
rect 735 45 737 47
rect 739 45 744 47
rect 746 45 757 47
rect 735 43 757 45
rect 761 47 767 49
rect 761 45 763 47
rect 765 45 767 47
rect 761 43 767 45
rect 775 46 777 59
rect 785 56 787 59
rect 781 54 787 56
rect 781 52 783 54
rect 785 52 787 54
rect 806 58 808 63
rect 816 58 818 63
rect 826 61 828 66
rect 781 50 787 52
rect 775 44 781 46
rect 633 40 642 42
rect 650 40 652 43
rect 657 40 659 43
rect 675 40 677 43
rect 685 40 687 43
rect 695 40 697 43
rect 717 40 719 43
rect 727 40 729 43
rect 737 40 739 43
rect 755 40 757 43
rect 762 40 764 43
rect 775 42 777 44
rect 779 42 781 44
rect 772 40 781 42
rect 640 37 642 40
rect 587 14 589 19
rect 597 14 599 19
rect 607 17 609 21
rect 518 8 520 12
rect 539 8 541 12
rect 546 8 548 12
rect 640 19 642 24
rect 627 8 629 12
rect 650 10 652 15
rect 657 10 659 15
rect 772 37 774 40
rect 785 37 787 50
rect 806 42 808 52
rect 816 49 818 52
rect 826 49 828 52
rect 812 47 818 49
rect 812 45 814 47
rect 816 45 818 47
rect 812 43 818 45
rect 822 47 828 49
rect 822 45 824 47
rect 826 45 828 47
rect 822 43 828 45
rect 802 40 808 42
rect 802 38 804 40
rect 806 38 808 40
rect 772 19 774 24
rect 675 8 677 12
rect 685 8 687 12
rect 695 8 697 12
rect 717 8 719 12
rect 727 8 729 12
rect 737 8 739 12
rect 755 10 757 15
rect 762 10 764 15
rect 802 36 808 38
rect 806 33 808 36
rect 813 33 815 43
rect 826 40 828 43
rect 826 17 828 22
rect 785 8 787 12
rect 806 8 808 12
rect 813 8 815 12
rect 831 5 833 7
rect 439 0 441 4
rect 424 -25 430 -23
rect 424 -27 426 -25
rect 428 -27 430 -25
rect 475 0 477 4
rect 495 0 497 4
rect 455 -9 457 -5
rect 465 -9 467 -5
rect 518 -3 520 2
rect 525 -3 527 2
rect 543 0 545 4
rect 553 0 555 4
rect 563 0 565 4
rect 585 0 587 4
rect 595 0 597 4
rect 605 0 607 4
rect 508 -12 510 -7
rect 424 -29 430 -27
rect 428 -30 430 -29
rect 439 -30 441 -27
rect 455 -30 457 -27
rect 428 -32 441 -30
rect 447 -32 457 -30
rect 465 -31 467 -27
rect 475 -30 477 -27
rect 431 -40 433 -32
rect 447 -36 449 -32
rect 440 -38 449 -36
rect 461 -33 467 -31
rect 461 -35 463 -33
rect 465 -35 467 -33
rect 461 -37 467 -35
rect 471 -32 477 -30
rect 471 -34 473 -32
rect 475 -34 477 -32
rect 471 -36 477 -34
rect 440 -40 442 -38
rect 444 -40 449 -38
rect 440 -42 449 -40
rect 465 -40 467 -37
rect 447 -45 449 -42
rect 457 -45 459 -41
rect 465 -42 469 -40
rect 467 -45 469 -42
rect 474 -45 476 -36
rect 495 -38 497 -25
rect 508 -28 510 -25
rect 623 -3 625 2
rect 630 -3 632 2
rect 653 0 655 4
rect 674 0 676 4
rect 681 0 683 4
rect 640 -12 642 -7
rect 727 0 729 4
rect 734 0 736 4
rect 744 0 746 4
rect 751 0 753 4
rect 761 0 763 4
rect 791 0 793 4
rect 798 0 800 4
rect 808 0 810 4
rect 815 0 817 4
rect 825 0 827 4
rect 694 -10 696 -5
rect 674 -24 676 -21
rect 640 -28 642 -25
rect 501 -30 510 -28
rect 501 -32 503 -30
rect 505 -32 507 -30
rect 518 -31 520 -28
rect 525 -31 527 -28
rect 543 -31 545 -28
rect 553 -31 555 -28
rect 563 -31 565 -28
rect 585 -31 587 -28
rect 595 -31 597 -28
rect 605 -31 607 -28
rect 623 -31 625 -28
rect 630 -31 632 -28
rect 640 -30 649 -28
rect 501 -34 507 -32
rect 495 -40 501 -38
rect 495 -42 497 -40
rect 499 -42 501 -40
rect 495 -44 501 -42
rect 431 -52 433 -49
rect 431 -54 436 -52
rect 434 -62 436 -54
rect 447 -58 449 -54
rect 457 -62 459 -54
rect 495 -47 497 -44
rect 505 -47 507 -34
rect 515 -33 521 -31
rect 515 -35 517 -33
rect 519 -35 521 -33
rect 515 -37 521 -35
rect 525 -33 547 -31
rect 525 -35 536 -33
rect 538 -35 543 -33
rect 545 -35 547 -33
rect 525 -37 547 -35
rect 551 -33 557 -31
rect 551 -35 553 -33
rect 555 -35 557 -33
rect 551 -37 557 -35
rect 561 -33 567 -31
rect 561 -35 563 -33
rect 565 -35 567 -33
rect 561 -37 567 -35
rect 583 -33 589 -31
rect 583 -35 585 -33
rect 587 -35 589 -33
rect 583 -37 589 -35
rect 593 -33 599 -31
rect 593 -35 595 -33
rect 597 -35 599 -33
rect 593 -37 599 -35
rect 603 -33 625 -31
rect 603 -35 605 -33
rect 607 -35 612 -33
rect 614 -35 625 -33
rect 603 -37 625 -35
rect 629 -33 635 -31
rect 629 -35 631 -33
rect 633 -35 635 -33
rect 629 -37 635 -35
rect 515 -40 517 -37
rect 525 -40 527 -37
rect 545 -40 547 -37
rect 552 -40 554 -37
rect 467 -62 469 -57
rect 474 -62 476 -57
rect 434 -64 459 -62
rect 495 -64 497 -60
rect 505 -62 507 -57
rect 515 -59 517 -54
rect 525 -59 527 -54
rect 563 -46 565 -37
rect 585 -46 587 -37
rect 596 -40 598 -37
rect 603 -40 605 -37
rect 623 -40 625 -37
rect 633 -40 635 -37
rect 643 -32 645 -30
rect 647 -32 649 -30
rect 643 -34 649 -32
rect 643 -47 645 -34
rect 653 -38 655 -25
rect 670 -26 676 -24
rect 670 -28 672 -26
rect 674 -28 676 -26
rect 670 -30 676 -28
rect 649 -40 655 -38
rect 674 -40 676 -30
rect 681 -31 683 -21
rect 710 -13 716 -11
rect 710 -15 712 -13
rect 714 -15 716 -13
rect 710 -17 719 -15
rect 717 -20 719 -17
rect 694 -31 696 -28
rect 680 -33 686 -31
rect 680 -35 682 -33
rect 684 -35 686 -33
rect 680 -37 686 -35
rect 690 -33 696 -31
rect 690 -35 692 -33
rect 694 -35 696 -33
rect 690 -37 696 -35
rect 684 -40 686 -37
rect 694 -40 696 -37
rect 649 -42 651 -40
rect 653 -42 655 -40
rect 649 -44 655 -42
rect 653 -47 655 -44
rect 623 -59 625 -54
rect 633 -59 635 -54
rect 545 -64 547 -60
rect 552 -64 554 -60
rect 563 -64 565 -60
rect 585 -64 587 -60
rect 596 -64 598 -60
rect 603 -64 605 -60
rect 643 -62 645 -57
rect 674 -51 676 -46
rect 684 -51 686 -46
rect 717 -46 719 -28
rect 727 -31 729 -16
rect 734 -21 736 -16
rect 733 -23 739 -21
rect 733 -25 735 -23
rect 737 -25 739 -23
rect 733 -27 739 -25
rect 744 -31 746 -16
rect 751 -26 753 -16
rect 774 -13 780 -11
rect 774 -15 776 -13
rect 778 -15 780 -13
rect 774 -17 783 -15
rect 723 -33 729 -31
rect 723 -35 725 -33
rect 727 -35 729 -33
rect 723 -37 729 -35
rect 727 -46 729 -37
rect 734 -33 746 -31
rect 750 -28 756 -26
rect 750 -30 752 -28
rect 754 -30 756 -28
rect 750 -32 756 -30
rect 734 -46 736 -33
rect 740 -39 746 -37
rect 740 -41 742 -39
rect 744 -41 746 -39
rect 740 -43 746 -41
rect 744 -46 746 -43
rect 751 -46 753 -32
rect 761 -36 763 -18
rect 781 -20 783 -17
rect 758 -38 764 -36
rect 758 -40 760 -38
rect 762 -40 764 -38
rect 758 -42 764 -40
rect 761 -45 763 -42
rect 694 -54 696 -49
rect 653 -64 655 -60
rect 717 -62 719 -52
rect 781 -46 783 -28
rect 791 -31 793 -16
rect 798 -21 800 -16
rect 797 -23 803 -21
rect 797 -25 799 -23
rect 801 -25 803 -23
rect 797 -27 803 -25
rect 808 -31 810 -16
rect 815 -26 817 -16
rect 787 -33 793 -31
rect 787 -35 789 -33
rect 791 -35 793 -33
rect 787 -37 793 -35
rect 791 -46 793 -37
rect 798 -33 810 -31
rect 814 -28 820 -26
rect 814 -30 816 -28
rect 818 -30 820 -28
rect 814 -32 820 -30
rect 798 -46 800 -33
rect 804 -39 810 -37
rect 804 -41 806 -39
rect 808 -41 810 -39
rect 804 -43 810 -41
rect 808 -46 810 -43
rect 815 -46 817 -32
rect 825 -36 827 -18
rect 822 -38 828 -36
rect 822 -40 824 -38
rect 826 -40 828 -38
rect 822 -42 828 -40
rect 825 -45 827 -42
rect 727 -58 729 -54
rect 734 -62 736 -54
rect 744 -59 746 -54
rect 751 -59 753 -54
rect 761 -59 763 -54
rect 717 -64 736 -62
rect 781 -62 783 -52
rect 791 -58 793 -54
rect 798 -62 800 -54
rect 808 -59 810 -54
rect 815 -59 817 -54
rect 825 -59 827 -54
rect 781 -64 800 -62
rect 434 -70 459 -68
rect 434 -78 436 -70
rect 447 -78 449 -74
rect 457 -78 459 -70
rect 467 -75 469 -70
rect 474 -75 476 -70
rect 495 -72 497 -68
rect 431 -80 436 -78
rect 431 -83 433 -80
rect 505 -75 507 -70
rect 545 -72 547 -68
rect 552 -72 554 -68
rect 563 -72 565 -68
rect 585 -72 587 -68
rect 596 -72 598 -68
rect 603 -72 605 -68
rect 515 -78 517 -73
rect 525 -78 527 -73
rect 447 -90 449 -87
rect 440 -92 449 -90
rect 457 -91 459 -87
rect 467 -90 469 -87
rect 431 -100 433 -92
rect 440 -94 442 -92
rect 444 -94 449 -92
rect 440 -96 449 -94
rect 465 -92 469 -90
rect 465 -95 467 -92
rect 447 -100 449 -96
rect 461 -97 467 -95
rect 474 -96 476 -87
rect 495 -88 497 -85
rect 495 -90 501 -88
rect 495 -92 497 -90
rect 499 -92 501 -90
rect 495 -94 501 -92
rect 461 -99 463 -97
rect 465 -99 467 -97
rect 428 -102 441 -100
rect 447 -102 457 -100
rect 461 -101 467 -99
rect 428 -103 430 -102
rect 424 -105 430 -103
rect 439 -105 441 -102
rect 455 -105 457 -102
rect 465 -105 467 -101
rect 471 -98 477 -96
rect 471 -100 473 -98
rect 475 -100 477 -98
rect 471 -102 477 -100
rect 475 -105 477 -102
rect 424 -107 426 -105
rect 428 -107 430 -105
rect 424 -109 430 -107
rect 455 -127 457 -123
rect 465 -127 467 -123
rect 439 -136 441 -132
rect 495 -107 497 -94
rect 505 -98 507 -85
rect 501 -100 507 -98
rect 501 -102 503 -100
rect 505 -102 507 -100
rect 515 -95 517 -92
rect 525 -95 527 -92
rect 545 -95 547 -92
rect 552 -95 554 -92
rect 563 -95 565 -86
rect 585 -95 587 -86
rect 623 -78 625 -73
rect 633 -78 635 -73
rect 643 -75 645 -70
rect 653 -72 655 -68
rect 717 -70 736 -68
rect 596 -95 598 -92
rect 603 -95 605 -92
rect 623 -95 625 -92
rect 633 -95 635 -92
rect 515 -97 521 -95
rect 515 -99 517 -97
rect 519 -99 521 -97
rect 515 -101 521 -99
rect 525 -97 547 -95
rect 525 -99 536 -97
rect 538 -99 543 -97
rect 545 -99 547 -97
rect 525 -101 547 -99
rect 551 -97 557 -95
rect 551 -99 553 -97
rect 555 -99 557 -97
rect 551 -101 557 -99
rect 561 -97 567 -95
rect 561 -99 563 -97
rect 565 -99 567 -97
rect 561 -101 567 -99
rect 583 -97 589 -95
rect 583 -99 585 -97
rect 587 -99 589 -97
rect 583 -101 589 -99
rect 593 -97 599 -95
rect 593 -99 595 -97
rect 597 -99 599 -97
rect 593 -101 599 -99
rect 603 -97 625 -95
rect 603 -99 605 -97
rect 607 -99 612 -97
rect 614 -99 625 -97
rect 603 -101 625 -99
rect 629 -97 635 -95
rect 629 -99 631 -97
rect 633 -99 635 -97
rect 629 -101 635 -99
rect 643 -98 645 -85
rect 653 -88 655 -85
rect 649 -90 655 -88
rect 649 -92 651 -90
rect 653 -92 655 -90
rect 674 -86 676 -81
rect 684 -86 686 -81
rect 694 -83 696 -78
rect 717 -80 719 -70
rect 727 -78 729 -74
rect 734 -78 736 -70
rect 781 -70 800 -68
rect 744 -78 746 -73
rect 751 -78 753 -73
rect 761 -78 763 -73
rect 649 -94 655 -92
rect 643 -100 649 -98
rect 501 -104 510 -102
rect 518 -104 520 -101
rect 525 -104 527 -101
rect 543 -104 545 -101
rect 553 -104 555 -101
rect 563 -104 565 -101
rect 585 -104 587 -101
rect 595 -104 597 -101
rect 605 -104 607 -101
rect 623 -104 625 -101
rect 630 -104 632 -101
rect 643 -102 645 -100
rect 647 -102 649 -100
rect 640 -104 649 -102
rect 508 -107 510 -104
rect 508 -125 510 -120
rect 475 -136 477 -132
rect 495 -136 497 -132
rect 518 -134 520 -129
rect 525 -134 527 -129
rect 640 -107 642 -104
rect 653 -107 655 -94
rect 674 -102 676 -92
rect 684 -95 686 -92
rect 694 -95 696 -92
rect 680 -97 686 -95
rect 680 -99 682 -97
rect 684 -99 686 -97
rect 680 -101 686 -99
rect 690 -97 696 -95
rect 690 -99 692 -97
rect 694 -99 696 -97
rect 690 -101 696 -99
rect 670 -104 676 -102
rect 670 -106 672 -104
rect 674 -106 676 -104
rect 640 -125 642 -120
rect 543 -136 545 -132
rect 553 -136 555 -132
rect 563 -136 565 -132
rect 585 -136 587 -132
rect 595 -136 597 -132
rect 605 -136 607 -132
rect 623 -134 625 -129
rect 630 -134 632 -129
rect 670 -108 676 -106
rect 674 -111 676 -108
rect 681 -111 683 -101
rect 694 -104 696 -101
rect 717 -104 719 -86
rect 727 -95 729 -86
rect 723 -97 729 -95
rect 723 -99 725 -97
rect 727 -99 729 -97
rect 723 -101 729 -99
rect 734 -99 736 -86
rect 744 -89 746 -86
rect 740 -91 746 -89
rect 740 -93 742 -91
rect 744 -93 746 -91
rect 740 -95 746 -93
rect 734 -101 746 -99
rect 751 -100 753 -86
rect 781 -80 783 -70
rect 791 -78 793 -74
rect 798 -78 800 -70
rect 808 -78 810 -73
rect 815 -78 817 -73
rect 825 -78 827 -73
rect 761 -90 763 -87
rect 758 -92 764 -90
rect 758 -94 760 -92
rect 762 -94 764 -92
rect 758 -96 764 -94
rect 717 -115 719 -112
rect 710 -117 719 -115
rect 727 -116 729 -101
rect 733 -107 739 -105
rect 733 -109 735 -107
rect 737 -109 739 -107
rect 733 -111 739 -109
rect 734 -116 736 -111
rect 744 -116 746 -101
rect 750 -102 756 -100
rect 750 -104 752 -102
rect 754 -104 756 -102
rect 750 -106 756 -104
rect 751 -116 753 -106
rect 761 -114 763 -96
rect 781 -104 783 -86
rect 791 -95 793 -86
rect 787 -97 793 -95
rect 787 -99 789 -97
rect 791 -99 793 -97
rect 787 -101 793 -99
rect 798 -99 800 -86
rect 808 -89 810 -86
rect 804 -91 810 -89
rect 804 -93 806 -91
rect 808 -93 810 -91
rect 804 -95 810 -93
rect 798 -101 810 -99
rect 815 -100 817 -86
rect 825 -90 827 -87
rect 822 -92 828 -90
rect 822 -94 824 -92
rect 826 -94 828 -92
rect 822 -96 828 -94
rect 710 -119 712 -117
rect 714 -119 716 -117
rect 710 -121 716 -119
rect 694 -127 696 -122
rect 653 -136 655 -132
rect 674 -136 676 -132
rect 681 -136 683 -132
rect 781 -115 783 -112
rect 774 -117 783 -115
rect 791 -116 793 -101
rect 797 -107 803 -105
rect 797 -109 799 -107
rect 801 -109 803 -107
rect 797 -111 803 -109
rect 798 -116 800 -111
rect 808 -116 810 -101
rect 814 -102 820 -100
rect 814 -104 816 -102
rect 818 -104 820 -102
rect 814 -106 820 -104
rect 815 -116 817 -106
rect 825 -114 827 -96
rect 774 -119 776 -117
rect 778 -119 780 -117
rect 774 -121 780 -119
rect 727 -136 729 -132
rect 734 -136 736 -132
rect 744 -136 746 -132
rect 751 -136 753 -132
rect 761 -136 763 -132
rect 791 -136 793 -132
rect 798 -136 800 -132
rect 808 -136 810 -132
rect 815 -136 817 -132
rect 825 -136 827 -132
rect 439 -144 441 -140
rect 424 -169 430 -167
rect 424 -171 426 -169
rect 428 -171 430 -169
rect 475 -144 477 -140
rect 495 -144 497 -140
rect 455 -153 457 -149
rect 465 -153 467 -149
rect 518 -147 520 -142
rect 525 -147 527 -142
rect 543 -144 545 -140
rect 553 -144 555 -140
rect 563 -144 565 -140
rect 585 -144 587 -140
rect 595 -144 597 -140
rect 605 -144 607 -140
rect 508 -156 510 -151
rect 424 -173 430 -171
rect 428 -174 430 -173
rect 439 -174 441 -171
rect 455 -174 457 -171
rect 428 -176 441 -174
rect 447 -176 457 -174
rect 465 -175 467 -171
rect 475 -174 477 -171
rect 431 -184 433 -176
rect 447 -180 449 -176
rect 440 -182 449 -180
rect 461 -177 467 -175
rect 461 -179 463 -177
rect 465 -179 467 -177
rect 461 -181 467 -179
rect 471 -176 477 -174
rect 471 -178 473 -176
rect 475 -178 477 -176
rect 471 -180 477 -178
rect 440 -184 442 -182
rect 444 -184 449 -182
rect 440 -186 449 -184
rect 465 -184 467 -181
rect 447 -189 449 -186
rect 457 -189 459 -185
rect 465 -186 469 -184
rect 467 -189 469 -186
rect 474 -189 476 -180
rect 495 -182 497 -169
rect 508 -172 510 -169
rect 623 -147 625 -142
rect 630 -147 632 -142
rect 653 -144 655 -140
rect 674 -144 676 -140
rect 681 -144 683 -140
rect 640 -156 642 -151
rect 727 -144 729 -140
rect 734 -144 736 -140
rect 744 -144 746 -140
rect 751 -144 753 -140
rect 761 -144 763 -140
rect 791 -144 793 -140
rect 798 -144 800 -140
rect 808 -144 810 -140
rect 815 -144 817 -140
rect 825 -144 827 -140
rect 694 -154 696 -149
rect 674 -168 676 -165
rect 640 -172 642 -169
rect 501 -174 510 -172
rect 501 -176 503 -174
rect 505 -176 507 -174
rect 518 -175 520 -172
rect 525 -175 527 -172
rect 543 -175 545 -172
rect 553 -175 555 -172
rect 563 -175 565 -172
rect 585 -175 587 -172
rect 595 -175 597 -172
rect 605 -175 607 -172
rect 623 -175 625 -172
rect 630 -175 632 -172
rect 640 -174 649 -172
rect 501 -178 507 -176
rect 495 -184 501 -182
rect 495 -186 497 -184
rect 499 -186 501 -184
rect 495 -188 501 -186
rect 431 -196 433 -193
rect 431 -198 436 -196
rect 434 -206 436 -198
rect 447 -202 449 -198
rect 457 -206 459 -198
rect 495 -191 497 -188
rect 505 -191 507 -178
rect 515 -177 521 -175
rect 515 -179 517 -177
rect 519 -179 521 -177
rect 515 -181 521 -179
rect 525 -177 547 -175
rect 525 -179 536 -177
rect 538 -179 543 -177
rect 545 -179 547 -177
rect 525 -181 547 -179
rect 551 -177 557 -175
rect 551 -179 553 -177
rect 555 -179 557 -177
rect 551 -181 557 -179
rect 561 -177 567 -175
rect 561 -179 563 -177
rect 565 -179 567 -177
rect 561 -181 567 -179
rect 583 -177 589 -175
rect 583 -179 585 -177
rect 587 -179 589 -177
rect 583 -181 589 -179
rect 593 -177 599 -175
rect 593 -179 595 -177
rect 597 -179 599 -177
rect 593 -181 599 -179
rect 603 -177 625 -175
rect 603 -179 605 -177
rect 607 -179 612 -177
rect 614 -179 625 -177
rect 603 -181 625 -179
rect 629 -177 635 -175
rect 629 -179 631 -177
rect 633 -179 635 -177
rect 629 -181 635 -179
rect 515 -184 517 -181
rect 525 -184 527 -181
rect 545 -184 547 -181
rect 552 -184 554 -181
rect 467 -206 469 -201
rect 474 -206 476 -201
rect 434 -208 459 -206
rect 495 -208 497 -204
rect 505 -206 507 -201
rect 515 -203 517 -198
rect 525 -203 527 -198
rect 563 -190 565 -181
rect 585 -190 587 -181
rect 596 -184 598 -181
rect 603 -184 605 -181
rect 623 -184 625 -181
rect 633 -184 635 -181
rect 643 -176 645 -174
rect 647 -176 649 -174
rect 643 -178 649 -176
rect 643 -191 645 -178
rect 653 -182 655 -169
rect 670 -170 676 -168
rect 670 -172 672 -170
rect 674 -172 676 -170
rect 670 -174 676 -172
rect 649 -184 655 -182
rect 674 -184 676 -174
rect 681 -175 683 -165
rect 710 -157 716 -155
rect 710 -159 712 -157
rect 714 -159 716 -157
rect 710 -161 719 -159
rect 717 -164 719 -161
rect 694 -175 696 -172
rect 680 -177 686 -175
rect 680 -179 682 -177
rect 684 -179 686 -177
rect 680 -181 686 -179
rect 690 -177 696 -175
rect 690 -179 692 -177
rect 694 -179 696 -177
rect 690 -181 696 -179
rect 684 -184 686 -181
rect 694 -184 696 -181
rect 649 -186 651 -184
rect 653 -186 655 -184
rect 649 -188 655 -186
rect 653 -191 655 -188
rect 623 -203 625 -198
rect 633 -203 635 -198
rect 545 -208 547 -204
rect 552 -208 554 -204
rect 563 -208 565 -204
rect 585 -208 587 -204
rect 596 -208 598 -204
rect 603 -208 605 -204
rect 643 -206 645 -201
rect 674 -195 676 -190
rect 684 -195 686 -190
rect 717 -190 719 -172
rect 727 -175 729 -160
rect 734 -165 736 -160
rect 733 -167 739 -165
rect 733 -169 735 -167
rect 737 -169 739 -167
rect 733 -171 739 -169
rect 744 -175 746 -160
rect 751 -170 753 -160
rect 774 -157 780 -155
rect 774 -159 776 -157
rect 778 -159 780 -157
rect 774 -161 783 -159
rect 723 -177 729 -175
rect 723 -179 725 -177
rect 727 -179 729 -177
rect 723 -181 729 -179
rect 727 -190 729 -181
rect 734 -177 746 -175
rect 750 -172 756 -170
rect 750 -174 752 -172
rect 754 -174 756 -172
rect 750 -176 756 -174
rect 734 -190 736 -177
rect 740 -183 746 -181
rect 740 -185 742 -183
rect 744 -185 746 -183
rect 740 -187 746 -185
rect 744 -190 746 -187
rect 751 -190 753 -176
rect 761 -180 763 -162
rect 781 -164 783 -161
rect 758 -182 764 -180
rect 758 -184 760 -182
rect 762 -184 764 -182
rect 758 -186 764 -184
rect 761 -189 763 -186
rect 694 -198 696 -193
rect 653 -208 655 -204
rect 717 -206 719 -196
rect 781 -190 783 -172
rect 791 -175 793 -160
rect 798 -165 800 -160
rect 797 -167 803 -165
rect 797 -169 799 -167
rect 801 -169 803 -167
rect 797 -171 803 -169
rect 808 -175 810 -160
rect 815 -170 817 -160
rect 787 -177 793 -175
rect 787 -179 789 -177
rect 791 -179 793 -177
rect 787 -181 793 -179
rect 791 -190 793 -181
rect 798 -177 810 -175
rect 814 -172 820 -170
rect 814 -174 816 -172
rect 818 -174 820 -172
rect 814 -176 820 -174
rect 798 -190 800 -177
rect 804 -183 810 -181
rect 804 -185 806 -183
rect 808 -185 810 -183
rect 804 -187 810 -185
rect 808 -190 810 -187
rect 815 -190 817 -176
rect 825 -180 827 -162
rect 822 -182 828 -180
rect 822 -184 824 -182
rect 826 -184 828 -182
rect 822 -186 828 -184
rect 825 -189 827 -186
rect 727 -202 729 -198
rect 734 -206 736 -198
rect 744 -203 746 -198
rect 751 -203 753 -198
rect 761 -203 763 -198
rect 717 -208 736 -206
rect 781 -206 783 -196
rect 791 -202 793 -198
rect 798 -206 800 -198
rect 808 -203 810 -198
rect 815 -203 817 -198
rect 825 -203 827 -198
rect 781 -208 800 -206
rect 434 -214 459 -212
rect 434 -222 436 -214
rect 447 -222 449 -218
rect 457 -222 459 -214
rect 467 -219 469 -214
rect 474 -219 476 -214
rect 495 -216 497 -212
rect 431 -224 436 -222
rect 431 -227 433 -224
rect 505 -219 507 -214
rect 545 -216 547 -212
rect 552 -216 554 -212
rect 563 -216 565 -212
rect 585 -216 587 -212
rect 596 -216 598 -212
rect 603 -216 605 -212
rect 515 -222 517 -217
rect 525 -222 527 -217
rect 447 -234 449 -231
rect 440 -236 449 -234
rect 457 -235 459 -231
rect 467 -234 469 -231
rect 431 -244 433 -236
rect 440 -238 442 -236
rect 444 -238 449 -236
rect 440 -240 449 -238
rect 465 -236 469 -234
rect 465 -239 467 -236
rect 447 -244 449 -240
rect 461 -241 467 -239
rect 474 -240 476 -231
rect 495 -232 497 -229
rect 495 -234 501 -232
rect 495 -236 497 -234
rect 499 -236 501 -234
rect 495 -238 501 -236
rect 461 -243 463 -241
rect 465 -243 467 -241
rect 428 -246 441 -244
rect 447 -246 457 -244
rect 461 -245 467 -243
rect 428 -247 430 -246
rect 424 -249 430 -247
rect 439 -249 441 -246
rect 455 -249 457 -246
rect 465 -249 467 -245
rect 471 -242 477 -240
rect 471 -244 473 -242
rect 475 -244 477 -242
rect 471 -246 477 -244
rect 475 -249 477 -246
rect 424 -251 426 -249
rect 428 -251 430 -249
rect 424 -253 430 -251
rect 455 -271 457 -267
rect 465 -271 467 -267
rect 439 -280 441 -276
rect 495 -251 497 -238
rect 505 -242 507 -229
rect 501 -244 507 -242
rect 501 -246 503 -244
rect 505 -246 507 -244
rect 515 -239 517 -236
rect 525 -239 527 -236
rect 545 -239 547 -236
rect 552 -239 554 -236
rect 563 -239 565 -230
rect 585 -239 587 -230
rect 623 -222 625 -217
rect 633 -222 635 -217
rect 643 -219 645 -214
rect 653 -216 655 -212
rect 717 -214 736 -212
rect 596 -239 598 -236
rect 603 -239 605 -236
rect 623 -239 625 -236
rect 633 -239 635 -236
rect 515 -241 521 -239
rect 515 -243 517 -241
rect 519 -243 521 -241
rect 515 -245 521 -243
rect 525 -241 547 -239
rect 525 -243 536 -241
rect 538 -243 543 -241
rect 545 -243 547 -241
rect 525 -245 547 -243
rect 551 -241 557 -239
rect 551 -243 553 -241
rect 555 -243 557 -241
rect 551 -245 557 -243
rect 561 -241 567 -239
rect 561 -243 563 -241
rect 565 -243 567 -241
rect 561 -245 567 -243
rect 583 -241 589 -239
rect 583 -243 585 -241
rect 587 -243 589 -241
rect 583 -245 589 -243
rect 593 -241 599 -239
rect 593 -243 595 -241
rect 597 -243 599 -241
rect 593 -245 599 -243
rect 603 -241 625 -239
rect 603 -243 605 -241
rect 607 -243 612 -241
rect 614 -243 625 -241
rect 603 -245 625 -243
rect 629 -241 635 -239
rect 629 -243 631 -241
rect 633 -243 635 -241
rect 629 -245 635 -243
rect 643 -242 645 -229
rect 653 -232 655 -229
rect 649 -234 655 -232
rect 649 -236 651 -234
rect 653 -236 655 -234
rect 674 -230 676 -225
rect 684 -230 686 -225
rect 694 -227 696 -222
rect 717 -224 719 -214
rect 727 -222 729 -218
rect 734 -222 736 -214
rect 781 -214 800 -212
rect 744 -222 746 -217
rect 751 -222 753 -217
rect 761 -222 763 -217
rect 649 -238 655 -236
rect 643 -244 649 -242
rect 501 -248 510 -246
rect 518 -248 520 -245
rect 525 -248 527 -245
rect 543 -248 545 -245
rect 553 -248 555 -245
rect 563 -248 565 -245
rect 585 -248 587 -245
rect 595 -248 597 -245
rect 605 -248 607 -245
rect 623 -248 625 -245
rect 630 -248 632 -245
rect 643 -246 645 -244
rect 647 -246 649 -244
rect 640 -248 649 -246
rect 508 -251 510 -248
rect 508 -269 510 -264
rect 475 -280 477 -276
rect 495 -280 497 -276
rect 518 -278 520 -273
rect 525 -278 527 -273
rect 640 -251 642 -248
rect 653 -251 655 -238
rect 674 -246 676 -236
rect 684 -239 686 -236
rect 694 -239 696 -236
rect 680 -241 686 -239
rect 680 -243 682 -241
rect 684 -243 686 -241
rect 680 -245 686 -243
rect 690 -241 696 -239
rect 690 -243 692 -241
rect 694 -243 696 -241
rect 690 -245 696 -243
rect 670 -248 676 -246
rect 670 -250 672 -248
rect 674 -250 676 -248
rect 640 -269 642 -264
rect 531 -280 533 -278
rect 543 -280 545 -276
rect 553 -280 555 -276
rect 563 -280 565 -276
rect 585 -280 587 -276
rect 595 -280 597 -276
rect 605 -280 607 -276
rect 623 -278 625 -273
rect 630 -278 632 -273
rect 670 -252 676 -250
rect 674 -255 676 -252
rect 681 -255 683 -245
rect 694 -248 696 -245
rect 717 -248 719 -230
rect 727 -239 729 -230
rect 723 -241 729 -239
rect 723 -243 725 -241
rect 727 -243 729 -241
rect 723 -245 729 -243
rect 734 -243 736 -230
rect 744 -233 746 -230
rect 740 -235 746 -233
rect 740 -237 742 -235
rect 744 -237 746 -235
rect 740 -239 746 -237
rect 734 -245 746 -243
rect 751 -244 753 -230
rect 781 -224 783 -214
rect 791 -222 793 -218
rect 798 -222 800 -214
rect 808 -222 810 -217
rect 815 -222 817 -217
rect 825 -222 827 -217
rect 761 -234 763 -231
rect 758 -236 764 -234
rect 758 -238 760 -236
rect 762 -238 764 -236
rect 758 -240 764 -238
rect 717 -259 719 -256
rect 710 -261 719 -259
rect 727 -260 729 -245
rect 733 -251 739 -249
rect 733 -253 735 -251
rect 737 -253 739 -251
rect 733 -255 739 -253
rect 734 -260 736 -255
rect 744 -260 746 -245
rect 750 -246 756 -244
rect 750 -248 752 -246
rect 754 -248 756 -246
rect 750 -250 756 -248
rect 751 -260 753 -250
rect 761 -258 763 -240
rect 781 -248 783 -230
rect 791 -239 793 -230
rect 787 -241 793 -239
rect 787 -243 789 -241
rect 791 -243 793 -241
rect 787 -245 793 -243
rect 798 -243 800 -230
rect 808 -233 810 -230
rect 804 -235 810 -233
rect 804 -237 806 -235
rect 808 -237 810 -235
rect 804 -239 810 -237
rect 798 -245 810 -243
rect 815 -244 817 -230
rect 825 -234 827 -231
rect 822 -236 828 -234
rect 822 -238 824 -236
rect 826 -238 828 -236
rect 822 -240 828 -238
rect 710 -263 712 -261
rect 714 -263 716 -261
rect 710 -265 716 -263
rect 694 -271 696 -266
rect 614 -280 616 -278
rect 653 -280 655 -276
rect 674 -280 676 -276
rect 681 -280 683 -276
rect 781 -259 783 -256
rect 774 -261 783 -259
rect 791 -260 793 -245
rect 797 -251 803 -249
rect 797 -253 799 -251
rect 801 -253 803 -251
rect 797 -255 803 -253
rect 798 -260 800 -255
rect 808 -260 810 -245
rect 814 -246 820 -244
rect 814 -248 816 -246
rect 818 -248 820 -246
rect 814 -250 820 -248
rect 815 -260 817 -250
rect 825 -258 827 -240
rect 774 -263 776 -261
rect 778 -263 780 -261
rect 774 -265 780 -263
rect 711 -280 713 -278
rect 727 -280 729 -276
rect 734 -280 736 -276
rect 744 -280 746 -276
rect 751 -280 753 -276
rect 761 -280 763 -276
rect 775 -280 777 -278
rect 791 -280 793 -276
rect 798 -280 800 -276
rect 808 -280 810 -276
rect 815 -280 817 -276
rect 825 -280 827 -276
<< ndif >>
rect 8 241 13 246
rect 6 239 13 241
rect 6 237 8 239
rect 10 237 13 239
rect 6 235 13 237
rect 15 235 20 246
rect 22 237 33 246
rect 35 243 40 246
rect 35 241 42 243
rect 48 241 53 246
rect 35 239 38 241
rect 40 239 42 241
rect 35 237 42 239
rect 46 239 53 241
rect 46 237 48 239
rect 50 237 53 239
rect 22 235 31 237
rect 24 229 31 235
rect 46 235 53 237
rect 55 235 60 246
rect 62 237 73 246
rect 75 243 80 246
rect 75 241 82 243
rect 108 241 113 248
rect 75 239 78 241
rect 80 239 82 241
rect 75 237 82 239
rect 86 239 93 241
rect 86 237 88 239
rect 90 237 93 239
rect 62 235 71 237
rect 24 227 27 229
rect 29 227 31 229
rect 24 225 31 227
rect 64 229 71 235
rect 86 235 93 237
rect 64 227 67 229
rect 69 227 71 229
rect 64 225 71 227
rect 88 228 93 235
rect 95 235 103 241
rect 95 233 98 235
rect 100 233 103 235
rect 95 231 103 233
rect 105 238 113 241
rect 105 236 108 238
rect 110 236 113 238
rect 105 234 113 236
rect 115 246 123 248
rect 115 244 118 246
rect 120 244 123 246
rect 115 234 123 244
rect 125 246 132 248
rect 125 244 128 246
rect 130 244 132 246
rect 125 239 132 244
rect 138 241 143 248
rect 125 237 128 239
rect 130 237 132 239
rect 125 234 132 237
rect 136 239 143 241
rect 136 237 138 239
rect 140 237 143 239
rect 136 235 143 237
rect 105 231 110 234
rect 95 228 100 231
rect 138 228 143 235
rect 145 228 150 248
rect 152 242 159 248
rect 187 242 194 248
rect 152 232 161 242
rect 152 230 155 232
rect 157 230 161 232
rect 152 228 161 230
rect 163 239 170 242
rect 163 237 166 239
rect 168 237 170 239
rect 163 235 170 237
rect 176 239 183 242
rect 176 237 178 239
rect 180 237 183 239
rect 176 235 183 237
rect 163 228 168 235
rect 178 228 183 235
rect 185 232 194 242
rect 185 230 189 232
rect 191 230 194 232
rect 185 228 194 230
rect 196 228 201 248
rect 203 241 208 248
rect 214 246 221 248
rect 214 244 216 246
rect 218 244 221 246
rect 203 239 210 241
rect 203 237 206 239
rect 208 237 210 239
rect 203 235 210 237
rect 214 239 221 244
rect 214 237 216 239
rect 218 237 221 239
rect 203 228 208 235
rect 214 234 221 237
rect 223 246 231 248
rect 223 244 226 246
rect 228 244 231 246
rect 223 234 231 244
rect 233 241 238 248
rect 265 242 272 248
rect 274 246 282 248
rect 274 244 277 246
rect 279 244 282 246
rect 274 242 282 244
rect 284 242 292 248
rect 233 238 241 241
rect 233 236 236 238
rect 238 236 241 238
rect 233 234 241 236
rect 236 231 241 234
rect 243 235 251 241
rect 243 233 246 235
rect 248 233 251 235
rect 243 231 251 233
rect 246 228 251 231
rect 253 239 260 241
rect 253 237 256 239
rect 258 237 260 239
rect 253 235 260 237
rect 265 235 270 242
rect 286 239 292 242
rect 294 246 301 248
rect 294 244 297 246
rect 299 244 301 246
rect 294 242 301 244
rect 294 239 299 242
rect 315 241 320 246
rect 313 239 320 241
rect 286 235 290 239
rect 253 228 258 235
rect 265 233 271 235
rect 265 231 267 233
rect 269 231 271 233
rect 265 229 271 231
rect 284 233 290 235
rect 313 237 315 239
rect 317 237 320 239
rect 313 235 320 237
rect 322 235 327 246
rect 329 237 340 246
rect 342 243 347 246
rect 342 241 349 243
rect 375 241 380 248
rect 342 239 345 241
rect 347 239 349 241
rect 342 237 349 239
rect 353 239 360 241
rect 353 237 355 239
rect 357 237 360 239
rect 329 235 338 237
rect 284 231 286 233
rect 288 231 290 233
rect 284 229 290 231
rect 331 229 338 235
rect 353 235 360 237
rect 331 227 334 229
rect 336 227 338 229
rect 331 225 338 227
rect 355 228 360 235
rect 362 235 370 241
rect 362 233 365 235
rect 367 233 370 235
rect 362 231 370 233
rect 372 238 380 241
rect 372 236 375 238
rect 377 236 380 238
rect 372 234 380 236
rect 382 246 390 248
rect 382 244 385 246
rect 387 244 390 246
rect 382 234 390 244
rect 392 246 399 248
rect 392 244 395 246
rect 397 244 399 246
rect 392 239 399 244
rect 405 241 410 248
rect 392 237 395 239
rect 397 237 399 239
rect 392 234 399 237
rect 403 239 410 241
rect 403 237 405 239
rect 407 237 410 239
rect 403 235 410 237
rect 372 231 377 234
rect 362 228 367 231
rect 405 228 410 235
rect 412 228 417 248
rect 419 242 426 248
rect 454 242 461 248
rect 419 232 428 242
rect 419 230 422 232
rect 424 230 428 232
rect 419 228 428 230
rect 430 239 437 242
rect 430 237 433 239
rect 435 237 437 239
rect 430 235 437 237
rect 443 239 450 242
rect 443 237 445 239
rect 447 237 450 239
rect 443 235 450 237
rect 430 228 435 235
rect 445 228 450 235
rect 452 232 461 242
rect 452 230 456 232
rect 458 230 461 232
rect 452 228 461 230
rect 463 228 468 248
rect 470 241 475 248
rect 481 246 488 248
rect 481 244 483 246
rect 485 244 488 246
rect 470 239 477 241
rect 470 237 473 239
rect 475 237 477 239
rect 470 235 477 237
rect 481 239 488 244
rect 481 237 483 239
rect 485 237 488 239
rect 470 228 475 235
rect 481 234 488 237
rect 490 246 498 248
rect 490 244 493 246
rect 495 244 498 246
rect 490 234 498 244
rect 500 241 505 248
rect 532 242 539 248
rect 541 246 549 248
rect 541 244 544 246
rect 546 244 549 246
rect 541 242 549 244
rect 551 242 559 248
rect 500 238 508 241
rect 500 236 503 238
rect 505 236 508 238
rect 500 234 508 236
rect 503 231 508 234
rect 510 235 518 241
rect 510 233 513 235
rect 515 233 518 235
rect 510 231 518 233
rect 513 228 518 231
rect 520 239 527 241
rect 520 237 523 239
rect 525 237 527 239
rect 520 235 527 237
rect 532 235 537 242
rect 553 239 559 242
rect 561 246 568 248
rect 561 244 564 246
rect 566 244 568 246
rect 561 242 568 244
rect 561 239 566 242
rect 582 241 587 246
rect 580 239 587 241
rect 553 235 557 239
rect 520 228 525 235
rect 532 233 538 235
rect 532 231 534 233
rect 536 231 538 233
rect 532 229 538 231
rect 551 233 557 235
rect 580 237 582 239
rect 584 237 587 239
rect 580 235 587 237
rect 589 235 594 246
rect 596 237 607 246
rect 609 243 614 246
rect 609 241 616 243
rect 642 241 647 248
rect 609 239 612 241
rect 614 239 616 241
rect 609 237 616 239
rect 620 239 627 241
rect 620 237 622 239
rect 624 237 627 239
rect 596 235 605 237
rect 551 231 553 233
rect 555 231 557 233
rect 551 229 557 231
rect 598 229 605 235
rect 620 235 627 237
rect 598 227 601 229
rect 603 227 605 229
rect 598 225 605 227
rect 622 228 627 235
rect 629 235 637 241
rect 629 233 632 235
rect 634 233 637 235
rect 629 231 637 233
rect 639 238 647 241
rect 639 236 642 238
rect 644 236 647 238
rect 639 234 647 236
rect 649 246 657 248
rect 649 244 652 246
rect 654 244 657 246
rect 649 234 657 244
rect 659 246 666 248
rect 659 244 662 246
rect 664 244 666 246
rect 659 239 666 244
rect 672 241 677 248
rect 659 237 662 239
rect 664 237 666 239
rect 659 234 666 237
rect 670 239 677 241
rect 670 237 672 239
rect 674 237 677 239
rect 670 235 677 237
rect 639 231 644 234
rect 629 228 634 231
rect 672 228 677 235
rect 679 228 684 248
rect 686 242 693 248
rect 721 242 728 248
rect 686 232 695 242
rect 686 230 689 232
rect 691 230 695 232
rect 686 228 695 230
rect 697 239 704 242
rect 697 237 700 239
rect 702 237 704 239
rect 697 235 704 237
rect 710 239 717 242
rect 710 237 712 239
rect 714 237 717 239
rect 710 235 717 237
rect 697 228 702 235
rect 712 228 717 235
rect 719 232 728 242
rect 719 230 723 232
rect 725 230 728 232
rect 719 228 728 230
rect 730 228 735 248
rect 737 241 742 248
rect 748 246 755 248
rect 748 244 750 246
rect 752 244 755 246
rect 737 239 744 241
rect 737 237 740 239
rect 742 237 744 239
rect 737 235 744 237
rect 748 239 755 244
rect 748 237 750 239
rect 752 237 755 239
rect 737 228 742 235
rect 748 234 755 237
rect 757 246 765 248
rect 757 244 760 246
rect 762 244 765 246
rect 757 234 765 244
rect 767 241 772 248
rect 799 242 806 248
rect 808 246 816 248
rect 808 244 811 246
rect 813 244 816 246
rect 808 242 816 244
rect 818 242 826 248
rect 767 238 775 241
rect 767 236 770 238
rect 772 236 775 238
rect 767 234 775 236
rect 770 231 775 234
rect 777 235 785 241
rect 777 233 780 235
rect 782 233 785 235
rect 777 231 785 233
rect 780 228 785 231
rect 787 239 794 241
rect 787 237 790 239
rect 792 237 794 239
rect 787 235 794 237
rect 799 235 804 242
rect 820 239 826 242
rect 828 246 835 248
rect 828 244 831 246
rect 833 244 835 246
rect 828 242 835 244
rect 828 239 833 242
rect 820 235 824 239
rect 787 228 792 235
rect 799 233 805 235
rect 799 231 801 233
rect 803 231 805 233
rect 799 229 805 231
rect 818 233 824 235
rect 818 231 820 233
rect 822 231 824 233
rect 818 229 824 231
rect 24 217 31 219
rect 24 215 27 217
rect 29 215 31 217
rect 24 209 31 215
rect 64 217 71 219
rect 64 215 67 217
rect 69 215 71 217
rect 6 207 13 209
rect 6 205 8 207
rect 10 205 13 207
rect 6 203 13 205
rect 8 198 13 203
rect 15 198 20 209
rect 22 207 31 209
rect 64 209 71 215
rect 46 207 53 209
rect 22 198 33 207
rect 35 205 42 207
rect 35 203 38 205
rect 40 203 42 205
rect 46 205 48 207
rect 50 205 53 207
rect 46 203 53 205
rect 35 201 42 203
rect 35 198 40 201
rect 48 198 53 203
rect 55 198 60 209
rect 62 207 71 209
rect 88 209 93 216
rect 86 207 93 209
rect 62 198 73 207
rect 75 205 82 207
rect 75 203 78 205
rect 80 203 82 205
rect 86 205 88 207
rect 90 205 93 207
rect 86 203 93 205
rect 95 213 100 216
rect 95 211 103 213
rect 95 209 98 211
rect 100 209 103 211
rect 95 203 103 209
rect 105 210 110 213
rect 105 208 113 210
rect 105 206 108 208
rect 110 206 113 208
rect 105 203 113 206
rect 75 201 82 203
rect 75 198 80 201
rect 108 196 113 203
rect 115 200 123 210
rect 115 198 118 200
rect 120 198 123 200
rect 115 196 123 198
rect 125 207 132 210
rect 138 209 143 216
rect 125 205 128 207
rect 130 205 132 207
rect 125 200 132 205
rect 136 207 143 209
rect 136 205 138 207
rect 140 205 143 207
rect 136 203 143 205
rect 125 198 128 200
rect 130 198 132 200
rect 125 196 132 198
rect 138 196 143 203
rect 145 196 150 216
rect 152 214 161 216
rect 152 212 155 214
rect 157 212 161 214
rect 152 202 161 212
rect 163 209 168 216
rect 178 209 183 216
rect 163 207 170 209
rect 163 205 166 207
rect 168 205 170 207
rect 163 202 170 205
rect 176 207 183 209
rect 176 205 178 207
rect 180 205 183 207
rect 176 202 183 205
rect 185 214 194 216
rect 185 212 189 214
rect 191 212 194 214
rect 185 202 194 212
rect 152 196 159 202
rect 187 196 194 202
rect 196 196 201 216
rect 203 209 208 216
rect 246 213 251 216
rect 236 210 241 213
rect 203 207 210 209
rect 203 205 206 207
rect 208 205 210 207
rect 203 203 210 205
rect 214 207 221 210
rect 214 205 216 207
rect 218 205 221 207
rect 203 196 208 203
rect 214 200 221 205
rect 214 198 216 200
rect 218 198 221 200
rect 214 196 221 198
rect 223 200 231 210
rect 223 198 226 200
rect 228 198 231 200
rect 223 196 231 198
rect 233 208 241 210
rect 233 206 236 208
rect 238 206 241 208
rect 233 203 241 206
rect 243 211 251 213
rect 243 209 246 211
rect 248 209 251 211
rect 243 203 251 209
rect 253 209 258 216
rect 265 213 271 215
rect 265 211 267 213
rect 269 211 271 213
rect 265 209 271 211
rect 284 213 290 215
rect 331 217 338 219
rect 331 215 334 217
rect 336 215 338 217
rect 284 211 286 213
rect 288 211 290 213
rect 284 209 290 211
rect 253 207 260 209
rect 253 205 256 207
rect 258 205 260 207
rect 253 203 260 205
rect 233 196 238 203
rect 265 202 270 209
rect 286 205 290 209
rect 331 209 338 215
rect 313 207 320 209
rect 313 205 315 207
rect 317 205 320 207
rect 286 202 292 205
rect 265 196 272 202
rect 274 200 282 202
rect 274 198 277 200
rect 279 198 282 200
rect 274 196 282 198
rect 284 196 292 202
rect 294 202 299 205
rect 313 203 320 205
rect 294 200 301 202
rect 294 198 297 200
rect 299 198 301 200
rect 315 198 320 203
rect 322 198 327 209
rect 329 207 338 209
rect 355 209 360 216
rect 353 207 360 209
rect 329 198 340 207
rect 342 205 349 207
rect 342 203 345 205
rect 347 203 349 205
rect 353 205 355 207
rect 357 205 360 207
rect 353 203 360 205
rect 362 213 367 216
rect 362 211 370 213
rect 362 209 365 211
rect 367 209 370 211
rect 362 203 370 209
rect 372 210 377 213
rect 372 208 380 210
rect 372 206 375 208
rect 377 206 380 208
rect 372 203 380 206
rect 342 201 349 203
rect 342 198 347 201
rect 294 196 301 198
rect 375 196 380 203
rect 382 200 390 210
rect 382 198 385 200
rect 387 198 390 200
rect 382 196 390 198
rect 392 207 399 210
rect 405 209 410 216
rect 392 205 395 207
rect 397 205 399 207
rect 392 200 399 205
rect 403 207 410 209
rect 403 205 405 207
rect 407 205 410 207
rect 403 203 410 205
rect 392 198 395 200
rect 397 198 399 200
rect 392 196 399 198
rect 405 196 410 203
rect 412 196 417 216
rect 419 214 428 216
rect 419 212 422 214
rect 424 212 428 214
rect 419 202 428 212
rect 430 209 435 216
rect 445 209 450 216
rect 430 207 437 209
rect 430 205 433 207
rect 435 205 437 207
rect 430 202 437 205
rect 443 207 450 209
rect 443 205 445 207
rect 447 205 450 207
rect 443 202 450 205
rect 452 214 461 216
rect 452 212 456 214
rect 458 212 461 214
rect 452 202 461 212
rect 419 196 426 202
rect 454 196 461 202
rect 463 196 468 216
rect 470 209 475 216
rect 513 213 518 216
rect 503 210 508 213
rect 470 207 477 209
rect 470 205 473 207
rect 475 205 477 207
rect 470 203 477 205
rect 481 207 488 210
rect 481 205 483 207
rect 485 205 488 207
rect 470 196 475 203
rect 481 200 488 205
rect 481 198 483 200
rect 485 198 488 200
rect 481 196 488 198
rect 490 200 498 210
rect 490 198 493 200
rect 495 198 498 200
rect 490 196 498 198
rect 500 208 508 210
rect 500 206 503 208
rect 505 206 508 208
rect 500 203 508 206
rect 510 211 518 213
rect 510 209 513 211
rect 515 209 518 211
rect 510 203 518 209
rect 520 209 525 216
rect 532 213 538 215
rect 532 211 534 213
rect 536 211 538 213
rect 532 209 538 211
rect 551 213 557 215
rect 598 217 605 219
rect 598 215 601 217
rect 603 215 605 217
rect 551 211 553 213
rect 555 211 557 213
rect 551 209 557 211
rect 520 207 527 209
rect 520 205 523 207
rect 525 205 527 207
rect 520 203 527 205
rect 500 196 505 203
rect 532 202 537 209
rect 553 205 557 209
rect 598 209 605 215
rect 580 207 587 209
rect 580 205 582 207
rect 584 205 587 207
rect 553 202 559 205
rect 532 196 539 202
rect 541 200 549 202
rect 541 198 544 200
rect 546 198 549 200
rect 541 196 549 198
rect 551 196 559 202
rect 561 202 566 205
rect 580 203 587 205
rect 561 200 568 202
rect 561 198 564 200
rect 566 198 568 200
rect 582 198 587 203
rect 589 198 594 209
rect 596 207 605 209
rect 622 209 627 216
rect 620 207 627 209
rect 596 198 607 207
rect 609 205 616 207
rect 609 203 612 205
rect 614 203 616 205
rect 620 205 622 207
rect 624 205 627 207
rect 620 203 627 205
rect 629 213 634 216
rect 629 211 637 213
rect 629 209 632 211
rect 634 209 637 211
rect 629 203 637 209
rect 639 210 644 213
rect 639 208 647 210
rect 639 206 642 208
rect 644 206 647 208
rect 639 203 647 206
rect 609 201 616 203
rect 609 198 614 201
rect 561 196 568 198
rect 642 196 647 203
rect 649 200 657 210
rect 649 198 652 200
rect 654 198 657 200
rect 649 196 657 198
rect 659 207 666 210
rect 672 209 677 216
rect 659 205 662 207
rect 664 205 666 207
rect 659 200 666 205
rect 670 207 677 209
rect 670 205 672 207
rect 674 205 677 207
rect 670 203 677 205
rect 659 198 662 200
rect 664 198 666 200
rect 659 196 666 198
rect 672 196 677 203
rect 679 196 684 216
rect 686 214 695 216
rect 686 212 689 214
rect 691 212 695 214
rect 686 202 695 212
rect 697 209 702 216
rect 712 209 717 216
rect 697 207 704 209
rect 697 205 700 207
rect 702 205 704 207
rect 697 202 704 205
rect 710 207 717 209
rect 710 205 712 207
rect 714 205 717 207
rect 710 202 717 205
rect 719 214 728 216
rect 719 212 723 214
rect 725 212 728 214
rect 719 202 728 212
rect 686 196 693 202
rect 721 196 728 202
rect 730 196 735 216
rect 737 209 742 216
rect 780 213 785 216
rect 770 210 775 213
rect 737 207 744 209
rect 737 205 740 207
rect 742 205 744 207
rect 737 203 744 205
rect 748 207 755 210
rect 748 205 750 207
rect 752 205 755 207
rect 737 196 742 203
rect 748 200 755 205
rect 748 198 750 200
rect 752 198 755 200
rect 748 196 755 198
rect 757 200 765 210
rect 757 198 760 200
rect 762 198 765 200
rect 757 196 765 198
rect 767 208 775 210
rect 767 206 770 208
rect 772 206 775 208
rect 767 203 775 206
rect 777 211 785 213
rect 777 209 780 211
rect 782 209 785 211
rect 777 203 785 209
rect 787 209 792 216
rect 799 213 805 215
rect 799 211 801 213
rect 803 211 805 213
rect 799 209 805 211
rect 818 213 824 215
rect 818 211 820 213
rect 822 211 824 213
rect 818 209 824 211
rect 787 207 794 209
rect 787 205 790 207
rect 792 205 794 207
rect 787 203 794 205
rect 767 196 772 203
rect 799 202 804 209
rect 820 205 824 209
rect 820 202 826 205
rect 799 196 806 202
rect 808 200 816 202
rect 808 198 811 200
rect 813 198 816 200
rect 808 196 816 198
rect 818 196 826 202
rect 828 202 833 205
rect 828 200 835 202
rect 828 198 831 200
rect 833 198 835 200
rect 828 196 835 198
rect 8 97 13 102
rect 6 95 13 97
rect 6 93 8 95
rect 10 93 13 95
rect 6 91 13 93
rect 15 91 20 102
rect 22 93 33 102
rect 35 99 40 102
rect 35 97 42 99
rect 48 97 53 102
rect 35 95 38 97
rect 40 95 42 97
rect 35 93 42 95
rect 46 95 53 97
rect 46 93 48 95
rect 50 93 53 95
rect 22 91 31 93
rect 24 85 31 91
rect 46 91 53 93
rect 55 91 60 102
rect 62 93 73 102
rect 75 99 80 102
rect 75 97 82 99
rect 108 97 113 104
rect 75 95 78 97
rect 80 95 82 97
rect 75 93 82 95
rect 86 95 93 97
rect 86 93 88 95
rect 90 93 93 95
rect 62 91 71 93
rect 24 83 27 85
rect 29 83 31 85
rect 24 81 31 83
rect 64 85 71 91
rect 86 91 93 93
rect 64 83 67 85
rect 69 83 71 85
rect 64 81 71 83
rect 88 84 93 91
rect 95 91 103 97
rect 95 89 98 91
rect 100 89 103 91
rect 95 87 103 89
rect 105 94 113 97
rect 105 92 108 94
rect 110 92 113 94
rect 105 90 113 92
rect 115 102 123 104
rect 115 100 118 102
rect 120 100 123 102
rect 115 90 123 100
rect 125 102 132 104
rect 125 100 128 102
rect 130 100 132 102
rect 125 95 132 100
rect 138 97 143 104
rect 125 93 128 95
rect 130 93 132 95
rect 125 90 132 93
rect 136 95 143 97
rect 136 93 138 95
rect 140 93 143 95
rect 136 91 143 93
rect 105 87 110 90
rect 95 84 100 87
rect 138 84 143 91
rect 145 84 150 104
rect 152 98 159 104
rect 187 98 194 104
rect 152 88 161 98
rect 152 86 155 88
rect 157 86 161 88
rect 152 84 161 86
rect 163 95 170 98
rect 163 93 166 95
rect 168 93 170 95
rect 163 91 170 93
rect 176 95 183 98
rect 176 93 178 95
rect 180 93 183 95
rect 176 91 183 93
rect 163 84 168 91
rect 178 84 183 91
rect 185 88 194 98
rect 185 86 189 88
rect 191 86 194 88
rect 185 84 194 86
rect 196 84 201 104
rect 203 97 208 104
rect 214 102 221 104
rect 214 100 216 102
rect 218 100 221 102
rect 203 95 210 97
rect 203 93 206 95
rect 208 93 210 95
rect 203 91 210 93
rect 214 95 221 100
rect 214 93 216 95
rect 218 93 221 95
rect 203 84 208 91
rect 214 90 221 93
rect 223 102 231 104
rect 223 100 226 102
rect 228 100 231 102
rect 223 90 231 100
rect 233 97 238 104
rect 265 98 272 104
rect 274 102 282 104
rect 274 100 277 102
rect 279 100 282 102
rect 274 98 282 100
rect 284 98 292 104
rect 233 94 241 97
rect 233 92 236 94
rect 238 92 241 94
rect 233 90 241 92
rect 236 87 241 90
rect 243 91 251 97
rect 243 89 246 91
rect 248 89 251 91
rect 243 87 251 89
rect 246 84 251 87
rect 253 95 260 97
rect 253 93 256 95
rect 258 93 260 95
rect 253 91 260 93
rect 265 91 270 98
rect 286 95 292 98
rect 294 102 301 104
rect 294 100 297 102
rect 299 100 301 102
rect 294 98 301 100
rect 294 95 299 98
rect 315 97 320 102
rect 313 95 320 97
rect 286 91 290 95
rect 253 84 258 91
rect 265 89 271 91
rect 265 87 267 89
rect 269 87 271 89
rect 265 85 271 87
rect 284 89 290 91
rect 313 93 315 95
rect 317 93 320 95
rect 313 91 320 93
rect 322 91 327 102
rect 329 93 340 102
rect 342 99 347 102
rect 342 97 349 99
rect 375 97 380 104
rect 342 95 345 97
rect 347 95 349 97
rect 342 93 349 95
rect 353 95 360 97
rect 353 93 355 95
rect 357 93 360 95
rect 329 91 338 93
rect 284 87 286 89
rect 288 87 290 89
rect 284 85 290 87
rect 331 85 338 91
rect 353 91 360 93
rect 331 83 334 85
rect 336 83 338 85
rect 331 81 338 83
rect 355 84 360 91
rect 362 91 370 97
rect 362 89 365 91
rect 367 89 370 91
rect 362 87 370 89
rect 372 94 380 97
rect 372 92 375 94
rect 377 92 380 94
rect 372 90 380 92
rect 382 102 390 104
rect 382 100 385 102
rect 387 100 390 102
rect 382 90 390 100
rect 392 102 399 104
rect 392 100 395 102
rect 397 100 399 102
rect 392 95 399 100
rect 405 97 410 104
rect 392 93 395 95
rect 397 93 399 95
rect 392 90 399 93
rect 403 95 410 97
rect 403 93 405 95
rect 407 93 410 95
rect 403 91 410 93
rect 372 87 377 90
rect 362 84 367 87
rect 405 84 410 91
rect 412 84 417 104
rect 419 98 426 104
rect 454 98 461 104
rect 419 88 428 98
rect 419 86 422 88
rect 424 86 428 88
rect 419 84 428 86
rect 430 95 437 98
rect 430 93 433 95
rect 435 93 437 95
rect 430 91 437 93
rect 443 95 450 98
rect 443 93 445 95
rect 447 93 450 95
rect 443 91 450 93
rect 430 84 435 91
rect 445 84 450 91
rect 452 88 461 98
rect 452 86 456 88
rect 458 86 461 88
rect 452 84 461 86
rect 463 84 468 104
rect 470 97 475 104
rect 481 102 488 104
rect 481 100 483 102
rect 485 100 488 102
rect 470 95 477 97
rect 470 93 473 95
rect 475 93 477 95
rect 470 91 477 93
rect 481 95 488 100
rect 481 93 483 95
rect 485 93 488 95
rect 470 84 475 91
rect 481 90 488 93
rect 490 102 498 104
rect 490 100 493 102
rect 495 100 498 102
rect 490 90 498 100
rect 500 97 505 104
rect 532 98 539 104
rect 541 102 549 104
rect 541 100 544 102
rect 546 100 549 102
rect 541 98 549 100
rect 551 98 559 104
rect 500 94 508 97
rect 500 92 503 94
rect 505 92 508 94
rect 500 90 508 92
rect 503 87 508 90
rect 510 91 518 97
rect 510 89 513 91
rect 515 89 518 91
rect 510 87 518 89
rect 513 84 518 87
rect 520 95 527 97
rect 520 93 523 95
rect 525 93 527 95
rect 520 91 527 93
rect 532 91 537 98
rect 553 95 559 98
rect 561 102 568 104
rect 561 100 564 102
rect 566 100 568 102
rect 561 98 568 100
rect 561 95 566 98
rect 582 97 587 102
rect 580 95 587 97
rect 553 91 557 95
rect 520 84 525 91
rect 532 89 538 91
rect 532 87 534 89
rect 536 87 538 89
rect 532 85 538 87
rect 551 89 557 91
rect 580 93 582 95
rect 584 93 587 95
rect 580 91 587 93
rect 589 91 594 102
rect 596 93 607 102
rect 609 99 614 102
rect 609 97 616 99
rect 642 97 647 104
rect 609 95 612 97
rect 614 95 616 97
rect 609 93 616 95
rect 620 95 627 97
rect 620 93 622 95
rect 624 93 627 95
rect 596 91 605 93
rect 551 87 553 89
rect 555 87 557 89
rect 551 85 557 87
rect 598 85 605 91
rect 620 91 627 93
rect 598 83 601 85
rect 603 83 605 85
rect 598 81 605 83
rect 622 84 627 91
rect 629 91 637 97
rect 629 89 632 91
rect 634 89 637 91
rect 629 87 637 89
rect 639 94 647 97
rect 639 92 642 94
rect 644 92 647 94
rect 639 90 647 92
rect 649 102 657 104
rect 649 100 652 102
rect 654 100 657 102
rect 649 90 657 100
rect 659 102 666 104
rect 659 100 662 102
rect 664 100 666 102
rect 659 95 666 100
rect 672 97 677 104
rect 659 93 662 95
rect 664 93 666 95
rect 659 90 666 93
rect 670 95 677 97
rect 670 93 672 95
rect 674 93 677 95
rect 670 91 677 93
rect 639 87 644 90
rect 629 84 634 87
rect 672 84 677 91
rect 679 84 684 104
rect 686 98 693 104
rect 721 98 728 104
rect 686 88 695 98
rect 686 86 689 88
rect 691 86 695 88
rect 686 84 695 86
rect 697 95 704 98
rect 697 93 700 95
rect 702 93 704 95
rect 697 91 704 93
rect 710 95 717 98
rect 710 93 712 95
rect 714 93 717 95
rect 710 91 717 93
rect 697 84 702 91
rect 712 84 717 91
rect 719 88 728 98
rect 719 86 723 88
rect 725 86 728 88
rect 719 84 728 86
rect 730 84 735 104
rect 737 97 742 104
rect 748 102 755 104
rect 748 100 750 102
rect 752 100 755 102
rect 737 95 744 97
rect 737 93 740 95
rect 742 93 744 95
rect 737 91 744 93
rect 748 95 755 100
rect 748 93 750 95
rect 752 93 755 95
rect 737 84 742 91
rect 748 90 755 93
rect 757 102 765 104
rect 757 100 760 102
rect 762 100 765 102
rect 757 90 765 100
rect 767 97 772 104
rect 799 98 806 104
rect 808 102 816 104
rect 808 100 811 102
rect 813 100 816 102
rect 808 98 816 100
rect 818 98 826 104
rect 767 94 775 97
rect 767 92 770 94
rect 772 92 775 94
rect 767 90 775 92
rect 770 87 775 90
rect 777 91 785 97
rect 777 89 780 91
rect 782 89 785 91
rect 777 87 785 89
rect 780 84 785 87
rect 787 95 794 97
rect 787 93 790 95
rect 792 93 794 95
rect 787 91 794 93
rect 799 91 804 98
rect 820 95 826 98
rect 828 102 835 104
rect 828 100 831 102
rect 833 100 835 102
rect 828 98 835 100
rect 828 95 833 98
rect 820 91 824 95
rect 787 84 792 91
rect 799 89 805 91
rect 799 87 801 89
rect 803 87 805 89
rect 799 85 805 87
rect 818 89 824 91
rect 818 87 820 89
rect 822 87 824 89
rect 818 85 824 87
rect 24 73 31 75
rect 24 71 27 73
rect 29 71 31 73
rect 24 65 31 71
rect 64 73 71 75
rect 64 71 67 73
rect 69 71 71 73
rect 6 63 13 65
rect 6 61 8 63
rect 10 61 13 63
rect 6 59 13 61
rect 8 54 13 59
rect 15 54 20 65
rect 22 63 31 65
rect 64 65 71 71
rect 46 63 53 65
rect 22 54 33 63
rect 35 61 42 63
rect 35 59 38 61
rect 40 59 42 61
rect 46 61 48 63
rect 50 61 53 63
rect 46 59 53 61
rect 35 57 42 59
rect 35 54 40 57
rect 48 54 53 59
rect 55 54 60 65
rect 62 63 71 65
rect 88 65 93 72
rect 86 63 93 65
rect 62 54 73 63
rect 75 61 82 63
rect 75 59 78 61
rect 80 59 82 61
rect 86 61 88 63
rect 90 61 93 63
rect 86 59 93 61
rect 95 69 100 72
rect 95 67 103 69
rect 95 65 98 67
rect 100 65 103 67
rect 95 59 103 65
rect 105 66 110 69
rect 105 64 113 66
rect 105 62 108 64
rect 110 62 113 64
rect 105 59 113 62
rect 75 57 82 59
rect 75 54 80 57
rect 108 52 113 59
rect 115 56 123 66
rect 115 54 118 56
rect 120 54 123 56
rect 115 52 123 54
rect 125 63 132 66
rect 138 65 143 72
rect 125 61 128 63
rect 130 61 132 63
rect 125 56 132 61
rect 136 63 143 65
rect 136 61 138 63
rect 140 61 143 63
rect 136 59 143 61
rect 125 54 128 56
rect 130 54 132 56
rect 125 52 132 54
rect 138 52 143 59
rect 145 52 150 72
rect 152 70 161 72
rect 152 68 155 70
rect 157 68 161 70
rect 152 58 161 68
rect 163 65 168 72
rect 178 65 183 72
rect 163 63 170 65
rect 163 61 166 63
rect 168 61 170 63
rect 163 58 170 61
rect 176 63 183 65
rect 176 61 178 63
rect 180 61 183 63
rect 176 58 183 61
rect 185 70 194 72
rect 185 68 189 70
rect 191 68 194 70
rect 185 58 194 68
rect 152 52 159 58
rect 187 52 194 58
rect 196 52 201 72
rect 203 65 208 72
rect 246 69 251 72
rect 236 66 241 69
rect 203 63 210 65
rect 203 61 206 63
rect 208 61 210 63
rect 203 59 210 61
rect 214 63 221 66
rect 214 61 216 63
rect 218 61 221 63
rect 203 52 208 59
rect 214 56 221 61
rect 214 54 216 56
rect 218 54 221 56
rect 214 52 221 54
rect 223 56 231 66
rect 223 54 226 56
rect 228 54 231 56
rect 223 52 231 54
rect 233 64 241 66
rect 233 62 236 64
rect 238 62 241 64
rect 233 59 241 62
rect 243 67 251 69
rect 243 65 246 67
rect 248 65 251 67
rect 243 59 251 65
rect 253 65 258 72
rect 265 69 271 71
rect 265 67 267 69
rect 269 67 271 69
rect 265 65 271 67
rect 284 69 290 71
rect 331 73 338 75
rect 331 71 334 73
rect 336 71 338 73
rect 284 67 286 69
rect 288 67 290 69
rect 284 65 290 67
rect 253 63 260 65
rect 253 61 256 63
rect 258 61 260 63
rect 253 59 260 61
rect 233 52 238 59
rect 265 58 270 65
rect 286 61 290 65
rect 331 65 338 71
rect 313 63 320 65
rect 313 61 315 63
rect 317 61 320 63
rect 286 58 292 61
rect 265 52 272 58
rect 274 56 282 58
rect 274 54 277 56
rect 279 54 282 56
rect 274 52 282 54
rect 284 52 292 58
rect 294 58 299 61
rect 313 59 320 61
rect 294 56 301 58
rect 294 54 297 56
rect 299 54 301 56
rect 315 54 320 59
rect 322 54 327 65
rect 329 63 338 65
rect 355 65 360 72
rect 353 63 360 65
rect 329 54 340 63
rect 342 61 349 63
rect 342 59 345 61
rect 347 59 349 61
rect 353 61 355 63
rect 357 61 360 63
rect 353 59 360 61
rect 362 69 367 72
rect 362 67 370 69
rect 362 65 365 67
rect 367 65 370 67
rect 362 59 370 65
rect 372 66 377 69
rect 372 64 380 66
rect 372 62 375 64
rect 377 62 380 64
rect 372 59 380 62
rect 342 57 349 59
rect 342 54 347 57
rect 294 52 301 54
rect 375 52 380 59
rect 382 56 390 66
rect 382 54 385 56
rect 387 54 390 56
rect 382 52 390 54
rect 392 63 399 66
rect 405 65 410 72
rect 392 61 395 63
rect 397 61 399 63
rect 392 56 399 61
rect 403 63 410 65
rect 403 61 405 63
rect 407 61 410 63
rect 403 59 410 61
rect 392 54 395 56
rect 397 54 399 56
rect 392 52 399 54
rect 405 52 410 59
rect 412 52 417 72
rect 419 70 428 72
rect 419 68 422 70
rect 424 68 428 70
rect 419 58 428 68
rect 430 65 435 72
rect 445 65 450 72
rect 430 63 437 65
rect 430 61 433 63
rect 435 61 437 63
rect 430 58 437 61
rect 443 63 450 65
rect 443 61 445 63
rect 447 61 450 63
rect 443 58 450 61
rect 452 70 461 72
rect 452 68 456 70
rect 458 68 461 70
rect 452 58 461 68
rect 419 52 426 58
rect 454 52 461 58
rect 463 52 468 72
rect 470 65 475 72
rect 513 69 518 72
rect 503 66 508 69
rect 470 63 477 65
rect 470 61 473 63
rect 475 61 477 63
rect 470 59 477 61
rect 481 63 488 66
rect 481 61 483 63
rect 485 61 488 63
rect 470 52 475 59
rect 481 56 488 61
rect 481 54 483 56
rect 485 54 488 56
rect 481 52 488 54
rect 490 56 498 66
rect 490 54 493 56
rect 495 54 498 56
rect 490 52 498 54
rect 500 64 508 66
rect 500 62 503 64
rect 505 62 508 64
rect 500 59 508 62
rect 510 67 518 69
rect 510 65 513 67
rect 515 65 518 67
rect 510 59 518 65
rect 520 65 525 72
rect 532 69 538 71
rect 532 67 534 69
rect 536 67 538 69
rect 532 65 538 67
rect 551 69 557 71
rect 598 73 605 75
rect 598 71 601 73
rect 603 71 605 73
rect 551 67 553 69
rect 555 67 557 69
rect 551 65 557 67
rect 520 63 527 65
rect 520 61 523 63
rect 525 61 527 63
rect 520 59 527 61
rect 500 52 505 59
rect 532 58 537 65
rect 553 61 557 65
rect 598 65 605 71
rect 580 63 587 65
rect 580 61 582 63
rect 584 61 587 63
rect 553 58 559 61
rect 532 52 539 58
rect 541 56 549 58
rect 541 54 544 56
rect 546 54 549 56
rect 541 52 549 54
rect 551 52 559 58
rect 561 58 566 61
rect 580 59 587 61
rect 561 56 568 58
rect 561 54 564 56
rect 566 54 568 56
rect 582 54 587 59
rect 589 54 594 65
rect 596 63 605 65
rect 622 65 627 72
rect 620 63 627 65
rect 596 54 607 63
rect 609 61 616 63
rect 609 59 612 61
rect 614 59 616 61
rect 620 61 622 63
rect 624 61 627 63
rect 620 59 627 61
rect 629 69 634 72
rect 629 67 637 69
rect 629 65 632 67
rect 634 65 637 67
rect 629 59 637 65
rect 639 66 644 69
rect 639 64 647 66
rect 639 62 642 64
rect 644 62 647 64
rect 639 59 647 62
rect 609 57 616 59
rect 609 54 614 57
rect 561 52 568 54
rect 642 52 647 59
rect 649 56 657 66
rect 649 54 652 56
rect 654 54 657 56
rect 649 52 657 54
rect 659 63 666 66
rect 672 65 677 72
rect 659 61 662 63
rect 664 61 666 63
rect 659 56 666 61
rect 670 63 677 65
rect 670 61 672 63
rect 674 61 677 63
rect 670 59 677 61
rect 659 54 662 56
rect 664 54 666 56
rect 659 52 666 54
rect 672 52 677 59
rect 679 52 684 72
rect 686 70 695 72
rect 686 68 689 70
rect 691 68 695 70
rect 686 58 695 68
rect 697 65 702 72
rect 712 65 717 72
rect 697 63 704 65
rect 697 61 700 63
rect 702 61 704 63
rect 697 58 704 61
rect 710 63 717 65
rect 710 61 712 63
rect 714 61 717 63
rect 710 58 717 61
rect 719 70 728 72
rect 719 68 723 70
rect 725 68 728 70
rect 719 58 728 68
rect 686 52 693 58
rect 721 52 728 58
rect 730 52 735 72
rect 737 65 742 72
rect 780 69 785 72
rect 770 66 775 69
rect 737 63 744 65
rect 737 61 740 63
rect 742 61 744 63
rect 737 59 744 61
rect 748 63 755 66
rect 748 61 750 63
rect 752 61 755 63
rect 737 52 742 59
rect 748 56 755 61
rect 748 54 750 56
rect 752 54 755 56
rect 748 52 755 54
rect 757 56 765 66
rect 757 54 760 56
rect 762 54 765 56
rect 757 52 765 54
rect 767 64 775 66
rect 767 62 770 64
rect 772 62 775 64
rect 767 59 775 62
rect 777 67 785 69
rect 777 65 780 67
rect 782 65 785 67
rect 777 59 785 65
rect 787 65 792 72
rect 799 69 805 71
rect 799 67 801 69
rect 803 67 805 69
rect 799 65 805 67
rect 818 69 824 71
rect 818 67 820 69
rect 822 67 824 69
rect 818 65 824 67
rect 787 63 794 65
rect 787 61 790 63
rect 792 61 794 63
rect 787 59 794 61
rect 767 52 772 59
rect 799 58 804 65
rect 820 61 824 65
rect 820 58 826 61
rect 799 52 806 58
rect 808 56 816 58
rect 808 54 811 56
rect 813 54 816 56
rect 808 52 816 54
rect 818 52 826 58
rect 828 58 833 61
rect 828 56 835 58
rect 828 54 831 56
rect 833 54 835 56
rect 828 52 835 54
rect 424 -42 431 -40
rect 424 -44 426 -42
rect 428 -44 431 -42
rect 424 -46 431 -44
rect 426 -49 431 -46
rect 433 -45 438 -40
rect 433 -49 447 -45
rect 438 -50 447 -49
rect 438 -52 440 -50
rect 442 -52 447 -50
rect 438 -54 447 -52
rect 449 -47 457 -45
rect 449 -49 452 -47
rect 454 -49 457 -47
rect 449 -54 457 -49
rect 459 -49 467 -45
rect 459 -51 462 -49
rect 464 -51 467 -49
rect 459 -54 467 -51
rect 462 -57 467 -54
rect 469 -57 474 -45
rect 476 -57 484 -45
rect 510 -47 515 -40
rect 488 -49 495 -47
rect 488 -51 490 -49
rect 492 -51 495 -49
rect 488 -53 495 -51
rect 478 -59 484 -57
rect 478 -61 480 -59
rect 482 -61 484 -59
rect 490 -60 495 -53
rect 497 -53 505 -47
rect 497 -55 500 -53
rect 502 -55 505 -53
rect 497 -57 505 -55
rect 507 -50 515 -47
rect 507 -52 510 -50
rect 512 -52 515 -50
rect 507 -54 515 -52
rect 517 -42 525 -40
rect 517 -44 520 -42
rect 522 -44 525 -42
rect 517 -54 525 -44
rect 527 -42 534 -40
rect 527 -44 530 -42
rect 532 -44 534 -42
rect 527 -49 534 -44
rect 540 -47 545 -40
rect 527 -51 530 -49
rect 532 -51 534 -49
rect 527 -54 534 -51
rect 538 -49 545 -47
rect 538 -51 540 -49
rect 542 -51 545 -49
rect 538 -53 545 -51
rect 507 -57 512 -54
rect 497 -60 502 -57
rect 478 -63 484 -61
rect 540 -60 545 -53
rect 547 -60 552 -40
rect 554 -46 561 -40
rect 589 -46 596 -40
rect 554 -56 563 -46
rect 554 -58 557 -56
rect 559 -58 563 -56
rect 554 -60 563 -58
rect 565 -49 572 -46
rect 565 -51 568 -49
rect 570 -51 572 -49
rect 565 -53 572 -51
rect 578 -49 585 -46
rect 578 -51 580 -49
rect 582 -51 585 -49
rect 578 -53 585 -51
rect 565 -60 570 -53
rect 580 -60 585 -53
rect 587 -56 596 -46
rect 587 -58 591 -56
rect 593 -58 596 -56
rect 587 -60 596 -58
rect 598 -60 603 -40
rect 605 -47 610 -40
rect 616 -42 623 -40
rect 616 -44 618 -42
rect 620 -44 623 -42
rect 605 -49 612 -47
rect 605 -51 608 -49
rect 610 -51 612 -49
rect 605 -53 612 -51
rect 616 -49 623 -44
rect 616 -51 618 -49
rect 620 -51 623 -49
rect 605 -60 610 -53
rect 616 -54 623 -51
rect 625 -42 633 -40
rect 625 -44 628 -42
rect 630 -44 633 -42
rect 625 -54 633 -44
rect 635 -47 640 -40
rect 667 -46 674 -40
rect 676 -42 684 -40
rect 676 -44 679 -42
rect 681 -44 684 -42
rect 676 -46 684 -44
rect 686 -46 694 -40
rect 635 -50 643 -47
rect 635 -52 638 -50
rect 640 -52 643 -50
rect 635 -54 643 -52
rect 638 -57 643 -54
rect 645 -53 653 -47
rect 645 -55 648 -53
rect 650 -55 653 -53
rect 645 -57 653 -55
rect 648 -60 653 -57
rect 655 -49 662 -47
rect 655 -51 658 -49
rect 660 -51 662 -49
rect 655 -53 662 -51
rect 667 -53 672 -46
rect 688 -49 694 -46
rect 696 -42 703 -40
rect 696 -44 699 -42
rect 701 -44 703 -42
rect 696 -46 703 -44
rect 756 -46 761 -45
rect 696 -49 701 -46
rect 710 -48 717 -46
rect 688 -53 692 -49
rect 655 -60 660 -53
rect 667 -55 673 -53
rect 667 -57 669 -55
rect 671 -57 673 -55
rect 667 -59 673 -57
rect 686 -55 692 -53
rect 710 -50 712 -48
rect 714 -50 717 -48
rect 710 -52 717 -50
rect 719 -48 727 -46
rect 719 -50 722 -48
rect 724 -50 727 -48
rect 719 -52 727 -50
rect 686 -57 688 -55
rect 690 -57 692 -55
rect 686 -59 692 -57
rect 721 -54 727 -52
rect 729 -54 734 -46
rect 736 -50 744 -46
rect 736 -52 739 -50
rect 741 -52 744 -50
rect 736 -54 744 -52
rect 746 -54 751 -46
rect 753 -50 761 -46
rect 753 -52 756 -50
rect 758 -52 761 -50
rect 753 -54 761 -52
rect 763 -47 770 -45
rect 820 -46 825 -45
rect 763 -49 766 -47
rect 768 -49 770 -47
rect 763 -51 770 -49
rect 774 -48 781 -46
rect 774 -50 776 -48
rect 778 -50 781 -48
rect 763 -54 768 -51
rect 774 -52 781 -50
rect 783 -48 791 -46
rect 783 -50 786 -48
rect 788 -50 791 -48
rect 783 -52 791 -50
rect 785 -54 791 -52
rect 793 -54 798 -46
rect 800 -50 808 -46
rect 800 -52 803 -50
rect 805 -52 808 -50
rect 800 -54 808 -52
rect 810 -54 815 -46
rect 817 -50 825 -46
rect 817 -52 820 -50
rect 822 -52 825 -50
rect 817 -54 825 -52
rect 827 -47 834 -45
rect 827 -49 830 -47
rect 832 -49 834 -47
rect 827 -51 834 -49
rect 827 -54 832 -51
rect 478 -71 484 -69
rect 478 -73 480 -71
rect 482 -73 484 -71
rect 478 -75 484 -73
rect 462 -78 467 -75
rect 438 -80 447 -78
rect 438 -82 440 -80
rect 442 -82 447 -80
rect 438 -83 447 -82
rect 426 -86 431 -83
rect 424 -88 431 -86
rect 424 -90 426 -88
rect 428 -90 431 -88
rect 424 -92 431 -90
rect 433 -87 447 -83
rect 449 -83 457 -78
rect 449 -85 452 -83
rect 454 -85 457 -83
rect 449 -87 457 -85
rect 459 -81 467 -78
rect 459 -83 462 -81
rect 464 -83 467 -81
rect 459 -87 467 -83
rect 469 -87 474 -75
rect 476 -87 484 -75
rect 490 -79 495 -72
rect 488 -81 495 -79
rect 488 -83 490 -81
rect 492 -83 495 -81
rect 488 -85 495 -83
rect 497 -75 502 -72
rect 497 -77 505 -75
rect 497 -79 500 -77
rect 502 -79 505 -77
rect 497 -85 505 -79
rect 507 -78 512 -75
rect 507 -80 515 -78
rect 507 -82 510 -80
rect 512 -82 515 -80
rect 507 -85 515 -82
rect 433 -92 438 -87
rect 510 -92 515 -85
rect 517 -88 525 -78
rect 517 -90 520 -88
rect 522 -90 525 -88
rect 517 -92 525 -90
rect 527 -81 534 -78
rect 540 -79 545 -72
rect 527 -83 530 -81
rect 532 -83 534 -81
rect 527 -88 534 -83
rect 538 -81 545 -79
rect 538 -83 540 -81
rect 542 -83 545 -81
rect 538 -85 545 -83
rect 527 -90 530 -88
rect 532 -90 534 -88
rect 527 -92 534 -90
rect 540 -92 545 -85
rect 547 -92 552 -72
rect 554 -74 563 -72
rect 554 -76 557 -74
rect 559 -76 563 -74
rect 554 -86 563 -76
rect 565 -79 570 -72
rect 580 -79 585 -72
rect 565 -81 572 -79
rect 565 -83 568 -81
rect 570 -83 572 -81
rect 565 -86 572 -83
rect 578 -81 585 -79
rect 578 -83 580 -81
rect 582 -83 585 -81
rect 578 -86 585 -83
rect 587 -74 596 -72
rect 587 -76 591 -74
rect 593 -76 596 -74
rect 587 -86 596 -76
rect 554 -92 561 -86
rect 589 -92 596 -86
rect 598 -92 603 -72
rect 605 -79 610 -72
rect 648 -75 653 -72
rect 638 -78 643 -75
rect 605 -81 612 -79
rect 605 -83 608 -81
rect 610 -83 612 -81
rect 605 -85 612 -83
rect 616 -81 623 -78
rect 616 -83 618 -81
rect 620 -83 623 -81
rect 605 -92 610 -85
rect 616 -88 623 -83
rect 616 -90 618 -88
rect 620 -90 623 -88
rect 616 -92 623 -90
rect 625 -88 633 -78
rect 625 -90 628 -88
rect 630 -90 633 -88
rect 625 -92 633 -90
rect 635 -80 643 -78
rect 635 -82 638 -80
rect 640 -82 643 -80
rect 635 -85 643 -82
rect 645 -77 653 -75
rect 645 -79 648 -77
rect 650 -79 653 -77
rect 645 -85 653 -79
rect 655 -79 660 -72
rect 667 -75 673 -73
rect 667 -77 669 -75
rect 671 -77 673 -75
rect 667 -79 673 -77
rect 686 -75 692 -73
rect 686 -77 688 -75
rect 690 -77 692 -75
rect 686 -79 692 -77
rect 655 -81 662 -79
rect 655 -83 658 -81
rect 660 -83 662 -81
rect 655 -85 662 -83
rect 635 -92 640 -85
rect 667 -86 672 -79
rect 688 -83 692 -79
rect 721 -80 727 -78
rect 710 -82 717 -80
rect 688 -86 694 -83
rect 667 -92 674 -86
rect 676 -88 684 -86
rect 676 -90 679 -88
rect 681 -90 684 -88
rect 676 -92 684 -90
rect 686 -92 694 -86
rect 696 -86 701 -83
rect 710 -84 712 -82
rect 714 -84 717 -82
rect 710 -86 717 -84
rect 719 -82 727 -80
rect 719 -84 722 -82
rect 724 -84 727 -82
rect 719 -86 727 -84
rect 729 -86 734 -78
rect 736 -80 744 -78
rect 736 -82 739 -80
rect 741 -82 744 -80
rect 736 -86 744 -82
rect 746 -86 751 -78
rect 753 -80 761 -78
rect 753 -82 756 -80
rect 758 -82 761 -80
rect 753 -86 761 -82
rect 696 -88 703 -86
rect 696 -90 699 -88
rect 701 -90 703 -88
rect 696 -92 703 -90
rect 756 -87 761 -86
rect 763 -81 768 -78
rect 785 -80 791 -78
rect 763 -83 770 -81
rect 763 -85 766 -83
rect 768 -85 770 -83
rect 763 -87 770 -85
rect 774 -82 781 -80
rect 774 -84 776 -82
rect 778 -84 781 -82
rect 774 -86 781 -84
rect 783 -82 791 -80
rect 783 -84 786 -82
rect 788 -84 791 -82
rect 783 -86 791 -84
rect 793 -86 798 -78
rect 800 -80 808 -78
rect 800 -82 803 -80
rect 805 -82 808 -80
rect 800 -86 808 -82
rect 810 -86 815 -78
rect 817 -80 825 -78
rect 817 -82 820 -80
rect 822 -82 825 -80
rect 817 -86 825 -82
rect 820 -87 825 -86
rect 827 -81 832 -78
rect 827 -83 834 -81
rect 827 -85 830 -83
rect 832 -85 834 -83
rect 827 -87 834 -85
rect 424 -186 431 -184
rect 424 -188 426 -186
rect 428 -188 431 -186
rect 424 -190 431 -188
rect 426 -193 431 -190
rect 433 -189 438 -184
rect 433 -193 447 -189
rect 438 -194 447 -193
rect 438 -196 440 -194
rect 442 -196 447 -194
rect 438 -198 447 -196
rect 449 -191 457 -189
rect 449 -193 452 -191
rect 454 -193 457 -191
rect 449 -198 457 -193
rect 459 -193 467 -189
rect 459 -195 462 -193
rect 464 -195 467 -193
rect 459 -198 467 -195
rect 462 -201 467 -198
rect 469 -201 474 -189
rect 476 -201 484 -189
rect 510 -191 515 -184
rect 488 -193 495 -191
rect 488 -195 490 -193
rect 492 -195 495 -193
rect 488 -197 495 -195
rect 478 -203 484 -201
rect 478 -205 480 -203
rect 482 -205 484 -203
rect 490 -204 495 -197
rect 497 -197 505 -191
rect 497 -199 500 -197
rect 502 -199 505 -197
rect 497 -201 505 -199
rect 507 -194 515 -191
rect 507 -196 510 -194
rect 512 -196 515 -194
rect 507 -198 515 -196
rect 517 -186 525 -184
rect 517 -188 520 -186
rect 522 -188 525 -186
rect 517 -198 525 -188
rect 527 -186 534 -184
rect 527 -188 530 -186
rect 532 -188 534 -186
rect 527 -193 534 -188
rect 540 -191 545 -184
rect 527 -195 530 -193
rect 532 -195 534 -193
rect 527 -198 534 -195
rect 538 -193 545 -191
rect 538 -195 540 -193
rect 542 -195 545 -193
rect 538 -197 545 -195
rect 507 -201 512 -198
rect 497 -204 502 -201
rect 478 -207 484 -205
rect 540 -204 545 -197
rect 547 -204 552 -184
rect 554 -190 561 -184
rect 589 -190 596 -184
rect 554 -200 563 -190
rect 554 -202 557 -200
rect 559 -202 563 -200
rect 554 -204 563 -202
rect 565 -193 572 -190
rect 565 -195 568 -193
rect 570 -195 572 -193
rect 565 -197 572 -195
rect 578 -193 585 -190
rect 578 -195 580 -193
rect 582 -195 585 -193
rect 578 -197 585 -195
rect 565 -204 570 -197
rect 580 -204 585 -197
rect 587 -200 596 -190
rect 587 -202 591 -200
rect 593 -202 596 -200
rect 587 -204 596 -202
rect 598 -204 603 -184
rect 605 -191 610 -184
rect 616 -186 623 -184
rect 616 -188 618 -186
rect 620 -188 623 -186
rect 605 -193 612 -191
rect 605 -195 608 -193
rect 610 -195 612 -193
rect 605 -197 612 -195
rect 616 -193 623 -188
rect 616 -195 618 -193
rect 620 -195 623 -193
rect 605 -204 610 -197
rect 616 -198 623 -195
rect 625 -186 633 -184
rect 625 -188 628 -186
rect 630 -188 633 -186
rect 625 -198 633 -188
rect 635 -191 640 -184
rect 667 -190 674 -184
rect 676 -186 684 -184
rect 676 -188 679 -186
rect 681 -188 684 -186
rect 676 -190 684 -188
rect 686 -190 694 -184
rect 635 -194 643 -191
rect 635 -196 638 -194
rect 640 -196 643 -194
rect 635 -198 643 -196
rect 638 -201 643 -198
rect 645 -197 653 -191
rect 645 -199 648 -197
rect 650 -199 653 -197
rect 645 -201 653 -199
rect 648 -204 653 -201
rect 655 -193 662 -191
rect 655 -195 658 -193
rect 660 -195 662 -193
rect 655 -197 662 -195
rect 667 -197 672 -190
rect 688 -193 694 -190
rect 696 -186 703 -184
rect 696 -188 699 -186
rect 701 -188 703 -186
rect 696 -190 703 -188
rect 756 -190 761 -189
rect 696 -193 701 -190
rect 710 -192 717 -190
rect 688 -197 692 -193
rect 655 -204 660 -197
rect 667 -199 673 -197
rect 667 -201 669 -199
rect 671 -201 673 -199
rect 667 -203 673 -201
rect 686 -199 692 -197
rect 710 -194 712 -192
rect 714 -194 717 -192
rect 710 -196 717 -194
rect 719 -192 727 -190
rect 719 -194 722 -192
rect 724 -194 727 -192
rect 719 -196 727 -194
rect 686 -201 688 -199
rect 690 -201 692 -199
rect 686 -203 692 -201
rect 721 -198 727 -196
rect 729 -198 734 -190
rect 736 -194 744 -190
rect 736 -196 739 -194
rect 741 -196 744 -194
rect 736 -198 744 -196
rect 746 -198 751 -190
rect 753 -194 761 -190
rect 753 -196 756 -194
rect 758 -196 761 -194
rect 753 -198 761 -196
rect 763 -191 770 -189
rect 820 -190 825 -189
rect 763 -193 766 -191
rect 768 -193 770 -191
rect 763 -195 770 -193
rect 774 -192 781 -190
rect 774 -194 776 -192
rect 778 -194 781 -192
rect 763 -198 768 -195
rect 774 -196 781 -194
rect 783 -192 791 -190
rect 783 -194 786 -192
rect 788 -194 791 -192
rect 783 -196 791 -194
rect 785 -198 791 -196
rect 793 -198 798 -190
rect 800 -194 808 -190
rect 800 -196 803 -194
rect 805 -196 808 -194
rect 800 -198 808 -196
rect 810 -198 815 -190
rect 817 -194 825 -190
rect 817 -196 820 -194
rect 822 -196 825 -194
rect 817 -198 825 -196
rect 827 -191 834 -189
rect 827 -193 830 -191
rect 832 -193 834 -191
rect 827 -195 834 -193
rect 827 -198 832 -195
rect 478 -215 484 -213
rect 478 -217 480 -215
rect 482 -217 484 -215
rect 478 -219 484 -217
rect 462 -222 467 -219
rect 438 -224 447 -222
rect 438 -226 440 -224
rect 442 -226 447 -224
rect 438 -227 447 -226
rect 426 -230 431 -227
rect 424 -232 431 -230
rect 424 -234 426 -232
rect 428 -234 431 -232
rect 424 -236 431 -234
rect 433 -231 447 -227
rect 449 -227 457 -222
rect 449 -229 452 -227
rect 454 -229 457 -227
rect 449 -231 457 -229
rect 459 -225 467 -222
rect 459 -227 462 -225
rect 464 -227 467 -225
rect 459 -231 467 -227
rect 469 -231 474 -219
rect 476 -231 484 -219
rect 490 -223 495 -216
rect 488 -225 495 -223
rect 488 -227 490 -225
rect 492 -227 495 -225
rect 488 -229 495 -227
rect 497 -219 502 -216
rect 497 -221 505 -219
rect 497 -223 500 -221
rect 502 -223 505 -221
rect 497 -229 505 -223
rect 507 -222 512 -219
rect 507 -224 515 -222
rect 507 -226 510 -224
rect 512 -226 515 -224
rect 507 -229 515 -226
rect 433 -236 438 -231
rect 510 -236 515 -229
rect 517 -232 525 -222
rect 517 -234 520 -232
rect 522 -234 525 -232
rect 517 -236 525 -234
rect 527 -225 534 -222
rect 540 -223 545 -216
rect 527 -227 530 -225
rect 532 -227 534 -225
rect 527 -232 534 -227
rect 538 -225 545 -223
rect 538 -227 540 -225
rect 542 -227 545 -225
rect 538 -229 545 -227
rect 527 -234 530 -232
rect 532 -234 534 -232
rect 527 -236 534 -234
rect 540 -236 545 -229
rect 547 -236 552 -216
rect 554 -218 563 -216
rect 554 -220 557 -218
rect 559 -220 563 -218
rect 554 -230 563 -220
rect 565 -223 570 -216
rect 580 -223 585 -216
rect 565 -225 572 -223
rect 565 -227 568 -225
rect 570 -227 572 -225
rect 565 -230 572 -227
rect 578 -225 585 -223
rect 578 -227 580 -225
rect 582 -227 585 -225
rect 578 -230 585 -227
rect 587 -218 596 -216
rect 587 -220 591 -218
rect 593 -220 596 -218
rect 587 -230 596 -220
rect 554 -236 561 -230
rect 589 -236 596 -230
rect 598 -236 603 -216
rect 605 -223 610 -216
rect 648 -219 653 -216
rect 638 -222 643 -219
rect 605 -225 612 -223
rect 605 -227 608 -225
rect 610 -227 612 -225
rect 605 -229 612 -227
rect 616 -225 623 -222
rect 616 -227 618 -225
rect 620 -227 623 -225
rect 605 -236 610 -229
rect 616 -232 623 -227
rect 616 -234 618 -232
rect 620 -234 623 -232
rect 616 -236 623 -234
rect 625 -232 633 -222
rect 625 -234 628 -232
rect 630 -234 633 -232
rect 625 -236 633 -234
rect 635 -224 643 -222
rect 635 -226 638 -224
rect 640 -226 643 -224
rect 635 -229 643 -226
rect 645 -221 653 -219
rect 645 -223 648 -221
rect 650 -223 653 -221
rect 645 -229 653 -223
rect 655 -223 660 -216
rect 667 -219 673 -217
rect 667 -221 669 -219
rect 671 -221 673 -219
rect 667 -223 673 -221
rect 686 -219 692 -217
rect 686 -221 688 -219
rect 690 -221 692 -219
rect 686 -223 692 -221
rect 655 -225 662 -223
rect 655 -227 658 -225
rect 660 -227 662 -225
rect 655 -229 662 -227
rect 635 -236 640 -229
rect 667 -230 672 -223
rect 688 -227 692 -223
rect 721 -224 727 -222
rect 710 -226 717 -224
rect 688 -230 694 -227
rect 667 -236 674 -230
rect 676 -232 684 -230
rect 676 -234 679 -232
rect 681 -234 684 -232
rect 676 -236 684 -234
rect 686 -236 694 -230
rect 696 -230 701 -227
rect 710 -228 712 -226
rect 714 -228 717 -226
rect 710 -230 717 -228
rect 719 -226 727 -224
rect 719 -228 722 -226
rect 724 -228 727 -226
rect 719 -230 727 -228
rect 729 -230 734 -222
rect 736 -224 744 -222
rect 736 -226 739 -224
rect 741 -226 744 -224
rect 736 -230 744 -226
rect 746 -230 751 -222
rect 753 -224 761 -222
rect 753 -226 756 -224
rect 758 -226 761 -224
rect 753 -230 761 -226
rect 696 -232 703 -230
rect 696 -234 699 -232
rect 701 -234 703 -232
rect 696 -236 703 -234
rect 756 -231 761 -230
rect 763 -225 768 -222
rect 785 -224 791 -222
rect 763 -227 770 -225
rect 763 -229 766 -227
rect 768 -229 770 -227
rect 763 -231 770 -229
rect 774 -226 781 -224
rect 774 -228 776 -226
rect 778 -228 781 -226
rect 774 -230 781 -228
rect 783 -226 791 -224
rect 783 -228 786 -226
rect 788 -228 791 -226
rect 783 -230 791 -228
rect 793 -230 798 -222
rect 800 -224 808 -222
rect 800 -226 803 -224
rect 805 -226 808 -224
rect 800 -230 808 -226
rect 810 -230 815 -222
rect 817 -224 825 -222
rect 817 -226 820 -224
rect 822 -226 825 -224
rect 817 -230 825 -226
rect 820 -231 825 -230
rect 827 -225 832 -222
rect 827 -227 834 -225
rect 827 -229 830 -227
rect 832 -229 834 -227
rect 827 -231 834 -229
<< pdif >>
rect 6 279 13 281
rect 6 277 8 279
rect 10 277 13 279
rect 6 268 13 277
rect 15 279 23 281
rect 15 277 18 279
rect 20 277 23 279
rect 15 272 23 277
rect 15 270 18 272
rect 20 270 23 272
rect 15 268 23 270
rect 25 279 31 281
rect 46 279 53 281
rect 25 277 33 279
rect 25 275 28 277
rect 30 275 33 277
rect 25 268 33 275
rect 27 261 33 268
rect 35 274 40 279
rect 46 277 48 279
rect 50 277 53 279
rect 35 272 42 274
rect 35 270 38 272
rect 40 270 42 272
rect 35 265 42 270
rect 46 268 53 277
rect 55 279 63 281
rect 55 277 58 279
rect 60 277 63 279
rect 55 272 63 277
rect 55 270 58 272
rect 60 270 63 272
rect 55 268 63 270
rect 65 279 71 281
rect 65 277 73 279
rect 65 275 68 277
rect 70 275 73 277
rect 65 268 73 275
rect 35 263 38 265
rect 40 263 42 265
rect 35 261 42 263
rect 67 261 73 268
rect 75 274 80 279
rect 88 276 93 288
rect 86 274 93 276
rect 75 272 82 274
rect 75 270 78 272
rect 80 270 82 272
rect 75 265 82 270
rect 75 263 78 265
rect 80 263 82 265
rect 86 272 88 274
rect 90 272 93 274
rect 86 267 93 272
rect 86 265 88 267
rect 90 265 93 267
rect 86 263 93 265
rect 95 286 104 288
rect 95 284 99 286
rect 101 284 104 286
rect 127 286 141 288
rect 127 285 134 286
rect 95 276 104 284
rect 111 276 116 285
rect 95 263 106 276
rect 108 267 116 276
rect 108 265 111 267
rect 113 265 116 267
rect 108 263 116 265
rect 75 261 82 263
rect 111 260 116 263
rect 118 260 123 285
rect 125 284 134 285
rect 136 284 141 286
rect 125 279 141 284
rect 125 277 134 279
rect 136 277 141 279
rect 125 260 141 277
rect 143 278 151 288
rect 143 276 146 278
rect 148 276 151 278
rect 143 271 151 276
rect 143 269 146 271
rect 148 269 151 271
rect 143 260 151 269
rect 153 286 161 288
rect 153 284 156 286
rect 158 284 161 286
rect 153 279 161 284
rect 153 277 156 279
rect 158 277 161 279
rect 153 260 161 277
rect 163 273 168 288
rect 178 273 183 288
rect 163 271 170 273
rect 163 269 166 271
rect 168 269 170 271
rect 163 264 170 269
rect 163 262 166 264
rect 168 262 170 264
rect 163 260 170 262
rect 176 271 183 273
rect 176 269 178 271
rect 180 269 183 271
rect 176 264 183 269
rect 176 262 178 264
rect 180 262 183 264
rect 176 260 183 262
rect 185 286 193 288
rect 185 284 188 286
rect 190 284 193 286
rect 185 279 193 284
rect 185 277 188 279
rect 190 277 193 279
rect 185 260 193 277
rect 195 278 203 288
rect 195 276 198 278
rect 200 276 203 278
rect 195 271 203 276
rect 195 269 198 271
rect 200 269 203 271
rect 195 260 203 269
rect 205 286 219 288
rect 205 284 210 286
rect 212 285 219 286
rect 242 286 251 288
rect 212 284 221 285
rect 205 279 221 284
rect 205 277 210 279
rect 212 277 221 279
rect 205 260 221 277
rect 223 260 228 285
rect 230 276 235 285
rect 242 284 245 286
rect 247 284 251 286
rect 242 276 251 284
rect 230 267 238 276
rect 230 265 233 267
rect 235 265 238 267
rect 230 263 238 265
rect 240 263 251 276
rect 253 276 258 288
rect 267 281 272 288
rect 265 279 272 281
rect 265 277 267 279
rect 269 277 272 279
rect 253 274 260 276
rect 265 275 272 277
rect 253 272 256 274
rect 258 272 260 274
rect 253 267 260 272
rect 267 267 272 275
rect 274 267 279 288
rect 281 286 290 288
rect 281 284 286 286
rect 288 284 290 286
rect 281 278 290 284
rect 313 279 320 281
rect 281 267 292 278
rect 253 265 256 267
rect 258 265 260 267
rect 253 263 260 265
rect 230 260 235 263
rect 284 260 292 267
rect 294 276 301 278
rect 294 274 297 276
rect 299 274 301 276
rect 294 269 301 274
rect 294 267 297 269
rect 299 267 301 269
rect 313 277 315 279
rect 317 277 320 279
rect 313 268 320 277
rect 322 279 330 281
rect 322 277 325 279
rect 327 277 330 279
rect 322 272 330 277
rect 322 270 325 272
rect 327 270 330 272
rect 322 268 330 270
rect 332 279 338 281
rect 332 277 340 279
rect 332 275 335 277
rect 337 275 340 277
rect 332 268 340 275
rect 294 265 301 267
rect 294 260 299 265
rect 334 261 340 268
rect 342 274 347 279
rect 355 276 360 288
rect 353 274 360 276
rect 342 272 349 274
rect 342 270 345 272
rect 347 270 349 272
rect 342 265 349 270
rect 342 263 345 265
rect 347 263 349 265
rect 353 272 355 274
rect 357 272 360 274
rect 353 267 360 272
rect 353 265 355 267
rect 357 265 360 267
rect 353 263 360 265
rect 362 286 371 288
rect 362 284 366 286
rect 368 284 371 286
rect 394 286 408 288
rect 394 285 401 286
rect 362 276 371 284
rect 378 276 383 285
rect 362 263 373 276
rect 375 267 383 276
rect 375 265 378 267
rect 380 265 383 267
rect 375 263 383 265
rect 342 261 349 263
rect 378 260 383 263
rect 385 260 390 285
rect 392 284 401 285
rect 403 284 408 286
rect 392 279 408 284
rect 392 277 401 279
rect 403 277 408 279
rect 392 260 408 277
rect 410 278 418 288
rect 410 276 413 278
rect 415 276 418 278
rect 410 271 418 276
rect 410 269 413 271
rect 415 269 418 271
rect 410 260 418 269
rect 420 286 428 288
rect 420 284 423 286
rect 425 284 428 286
rect 420 279 428 284
rect 420 277 423 279
rect 425 277 428 279
rect 420 260 428 277
rect 430 273 435 288
rect 445 273 450 288
rect 430 271 437 273
rect 430 269 433 271
rect 435 269 437 271
rect 430 264 437 269
rect 430 262 433 264
rect 435 262 437 264
rect 430 260 437 262
rect 443 271 450 273
rect 443 269 445 271
rect 447 269 450 271
rect 443 264 450 269
rect 443 262 445 264
rect 447 262 450 264
rect 443 260 450 262
rect 452 286 460 288
rect 452 284 455 286
rect 457 284 460 286
rect 452 279 460 284
rect 452 277 455 279
rect 457 277 460 279
rect 452 260 460 277
rect 462 278 470 288
rect 462 276 465 278
rect 467 276 470 278
rect 462 271 470 276
rect 462 269 465 271
rect 467 269 470 271
rect 462 260 470 269
rect 472 286 486 288
rect 472 284 477 286
rect 479 285 486 286
rect 509 286 518 288
rect 479 284 488 285
rect 472 279 488 284
rect 472 277 477 279
rect 479 277 488 279
rect 472 260 488 277
rect 490 260 495 285
rect 497 276 502 285
rect 509 284 512 286
rect 514 284 518 286
rect 509 276 518 284
rect 497 267 505 276
rect 497 265 500 267
rect 502 265 505 267
rect 497 263 505 265
rect 507 263 518 276
rect 520 276 525 288
rect 534 281 539 288
rect 532 279 539 281
rect 532 277 534 279
rect 536 277 539 279
rect 520 274 527 276
rect 532 275 539 277
rect 520 272 523 274
rect 525 272 527 274
rect 520 267 527 272
rect 534 267 539 275
rect 541 267 546 288
rect 548 286 557 288
rect 548 284 553 286
rect 555 284 557 286
rect 548 278 557 284
rect 580 279 587 281
rect 548 267 559 278
rect 520 265 523 267
rect 525 265 527 267
rect 520 263 527 265
rect 497 260 502 263
rect 551 260 559 267
rect 561 276 568 278
rect 561 274 564 276
rect 566 274 568 276
rect 561 269 568 274
rect 561 267 564 269
rect 566 267 568 269
rect 580 277 582 279
rect 584 277 587 279
rect 580 268 587 277
rect 589 279 597 281
rect 589 277 592 279
rect 594 277 597 279
rect 589 272 597 277
rect 589 270 592 272
rect 594 270 597 272
rect 589 268 597 270
rect 599 279 605 281
rect 599 277 607 279
rect 599 275 602 277
rect 604 275 607 277
rect 599 268 607 275
rect 561 265 568 267
rect 561 260 566 265
rect 601 261 607 268
rect 609 274 614 279
rect 622 276 627 288
rect 620 274 627 276
rect 609 272 616 274
rect 609 270 612 272
rect 614 270 616 272
rect 609 265 616 270
rect 609 263 612 265
rect 614 263 616 265
rect 620 272 622 274
rect 624 272 627 274
rect 620 267 627 272
rect 620 265 622 267
rect 624 265 627 267
rect 620 263 627 265
rect 629 286 638 288
rect 629 284 633 286
rect 635 284 638 286
rect 661 286 675 288
rect 661 285 668 286
rect 629 276 638 284
rect 645 276 650 285
rect 629 263 640 276
rect 642 267 650 276
rect 642 265 645 267
rect 647 265 650 267
rect 642 263 650 265
rect 609 261 616 263
rect 645 260 650 263
rect 652 260 657 285
rect 659 284 668 285
rect 670 284 675 286
rect 659 279 675 284
rect 659 277 668 279
rect 670 277 675 279
rect 659 260 675 277
rect 677 278 685 288
rect 677 276 680 278
rect 682 276 685 278
rect 677 271 685 276
rect 677 269 680 271
rect 682 269 685 271
rect 677 260 685 269
rect 687 286 695 288
rect 687 284 690 286
rect 692 284 695 286
rect 687 279 695 284
rect 687 277 690 279
rect 692 277 695 279
rect 687 260 695 277
rect 697 273 702 288
rect 712 273 717 288
rect 697 271 704 273
rect 697 269 700 271
rect 702 269 704 271
rect 697 264 704 269
rect 697 262 700 264
rect 702 262 704 264
rect 697 260 704 262
rect 710 271 717 273
rect 710 269 712 271
rect 714 269 717 271
rect 710 264 717 269
rect 710 262 712 264
rect 714 262 717 264
rect 710 260 717 262
rect 719 286 727 288
rect 719 284 722 286
rect 724 284 727 286
rect 719 279 727 284
rect 719 277 722 279
rect 724 277 727 279
rect 719 260 727 277
rect 729 278 737 288
rect 729 276 732 278
rect 734 276 737 278
rect 729 271 737 276
rect 729 269 732 271
rect 734 269 737 271
rect 729 260 737 269
rect 739 286 753 288
rect 739 284 744 286
rect 746 285 753 286
rect 776 286 785 288
rect 746 284 755 285
rect 739 279 755 284
rect 739 277 744 279
rect 746 277 755 279
rect 739 260 755 277
rect 757 260 762 285
rect 764 276 769 285
rect 776 284 779 286
rect 781 284 785 286
rect 776 276 785 284
rect 764 267 772 276
rect 764 265 767 267
rect 769 265 772 267
rect 764 263 772 265
rect 774 263 785 276
rect 787 276 792 288
rect 801 281 806 288
rect 799 279 806 281
rect 799 277 801 279
rect 803 277 806 279
rect 787 274 794 276
rect 799 275 806 277
rect 787 272 790 274
rect 792 272 794 274
rect 787 267 794 272
rect 801 267 806 275
rect 808 267 813 288
rect 815 286 824 288
rect 815 284 820 286
rect 822 284 824 286
rect 815 278 824 284
rect 815 267 826 278
rect 787 265 790 267
rect 792 265 794 267
rect 787 263 794 265
rect 764 260 769 263
rect 818 260 826 267
rect 828 276 835 278
rect 828 274 831 276
rect 833 274 835 276
rect 828 269 835 274
rect 828 267 831 269
rect 833 267 835 269
rect 828 265 835 267
rect 828 260 833 265
rect 27 176 33 183
rect 6 167 13 176
rect 6 165 8 167
rect 10 165 13 167
rect 6 163 13 165
rect 15 174 23 176
rect 15 172 18 174
rect 20 172 23 174
rect 15 167 23 172
rect 15 165 18 167
rect 20 165 23 167
rect 15 163 23 165
rect 25 169 33 176
rect 25 167 28 169
rect 30 167 33 169
rect 25 165 33 167
rect 35 180 42 183
rect 35 178 38 180
rect 40 178 42 180
rect 35 172 42 178
rect 67 176 73 183
rect 35 170 38 172
rect 40 170 42 172
rect 35 168 42 170
rect 35 165 40 168
rect 46 167 53 176
rect 46 165 48 167
rect 50 165 53 167
rect 25 163 31 165
rect 46 163 53 165
rect 55 174 63 176
rect 55 172 58 174
rect 60 172 63 174
rect 55 167 63 172
rect 55 165 58 167
rect 60 165 63 167
rect 55 163 63 165
rect 65 169 73 176
rect 65 167 68 169
rect 70 167 73 169
rect 65 165 73 167
rect 75 181 82 183
rect 111 181 116 184
rect 75 179 78 181
rect 80 179 82 181
rect 75 174 82 179
rect 75 172 78 174
rect 80 172 82 174
rect 75 170 82 172
rect 86 179 93 181
rect 86 177 88 179
rect 90 177 93 179
rect 86 172 93 177
rect 86 170 88 172
rect 90 170 93 172
rect 75 165 80 170
rect 86 168 93 170
rect 65 163 71 165
rect 88 156 93 168
rect 95 168 106 181
rect 108 179 116 181
rect 108 177 111 179
rect 113 177 116 179
rect 108 168 116 177
rect 95 160 104 168
rect 95 158 99 160
rect 101 158 104 160
rect 111 159 116 168
rect 118 159 123 184
rect 125 167 141 184
rect 125 165 134 167
rect 136 165 141 167
rect 125 160 141 165
rect 125 159 134 160
rect 95 156 104 158
rect 127 158 134 159
rect 136 158 141 160
rect 127 156 141 158
rect 143 175 151 184
rect 143 173 146 175
rect 148 173 151 175
rect 143 168 151 173
rect 143 166 146 168
rect 148 166 151 168
rect 143 156 151 166
rect 153 167 161 184
rect 153 165 156 167
rect 158 165 161 167
rect 153 160 161 165
rect 153 158 156 160
rect 158 158 161 160
rect 153 156 161 158
rect 163 182 170 184
rect 163 180 166 182
rect 168 180 170 182
rect 163 175 170 180
rect 163 173 166 175
rect 168 173 170 175
rect 163 171 170 173
rect 176 182 183 184
rect 176 180 178 182
rect 180 180 183 182
rect 176 175 183 180
rect 176 173 178 175
rect 180 173 183 175
rect 176 171 183 173
rect 163 156 168 171
rect 178 156 183 171
rect 185 167 193 184
rect 185 165 188 167
rect 190 165 193 167
rect 185 160 193 165
rect 185 158 188 160
rect 190 158 193 160
rect 185 156 193 158
rect 195 175 203 184
rect 195 173 198 175
rect 200 173 203 175
rect 195 168 203 173
rect 195 166 198 168
rect 200 166 203 168
rect 195 156 203 166
rect 205 167 221 184
rect 205 165 210 167
rect 212 165 221 167
rect 205 160 221 165
rect 205 158 210 160
rect 212 159 221 160
rect 223 159 228 184
rect 230 181 235 184
rect 230 179 238 181
rect 230 177 233 179
rect 235 177 238 179
rect 230 168 238 177
rect 240 168 251 181
rect 230 159 235 168
rect 242 160 251 168
rect 212 158 219 159
rect 205 156 219 158
rect 242 158 245 160
rect 247 158 251 160
rect 242 156 251 158
rect 253 179 260 181
rect 253 177 256 179
rect 258 177 260 179
rect 284 177 292 184
rect 253 172 260 177
rect 253 170 256 172
rect 258 170 260 172
rect 253 168 260 170
rect 267 169 272 177
rect 253 156 258 168
rect 265 167 272 169
rect 265 165 267 167
rect 269 165 272 167
rect 265 163 272 165
rect 267 156 272 163
rect 274 156 279 177
rect 281 166 292 177
rect 294 179 299 184
rect 294 177 301 179
rect 294 175 297 177
rect 299 175 301 177
rect 334 176 340 183
rect 294 170 301 175
rect 294 168 297 170
rect 299 168 301 170
rect 294 166 301 168
rect 313 167 320 176
rect 281 160 290 166
rect 313 165 315 167
rect 317 165 320 167
rect 313 163 320 165
rect 322 174 330 176
rect 322 172 325 174
rect 327 172 330 174
rect 322 167 330 172
rect 322 165 325 167
rect 327 165 330 167
rect 322 163 330 165
rect 332 169 340 176
rect 332 167 335 169
rect 337 167 340 169
rect 332 165 340 167
rect 342 181 349 183
rect 378 181 383 184
rect 342 179 345 181
rect 347 179 349 181
rect 342 174 349 179
rect 342 172 345 174
rect 347 172 349 174
rect 342 170 349 172
rect 353 179 360 181
rect 353 177 355 179
rect 357 177 360 179
rect 353 172 360 177
rect 353 170 355 172
rect 357 170 360 172
rect 342 165 347 170
rect 353 168 360 170
rect 332 163 338 165
rect 281 158 286 160
rect 288 158 290 160
rect 281 156 290 158
rect 355 156 360 168
rect 362 168 373 181
rect 375 179 383 181
rect 375 177 378 179
rect 380 177 383 179
rect 375 168 383 177
rect 362 160 371 168
rect 362 158 366 160
rect 368 158 371 160
rect 378 159 383 168
rect 385 159 390 184
rect 392 167 408 184
rect 392 165 401 167
rect 403 165 408 167
rect 392 160 408 165
rect 392 159 401 160
rect 362 156 371 158
rect 394 158 401 159
rect 403 158 408 160
rect 394 156 408 158
rect 410 175 418 184
rect 410 173 413 175
rect 415 173 418 175
rect 410 168 418 173
rect 410 166 413 168
rect 415 166 418 168
rect 410 156 418 166
rect 420 167 428 184
rect 420 165 423 167
rect 425 165 428 167
rect 420 160 428 165
rect 420 158 423 160
rect 425 158 428 160
rect 420 156 428 158
rect 430 182 437 184
rect 430 180 433 182
rect 435 180 437 182
rect 430 175 437 180
rect 430 173 433 175
rect 435 173 437 175
rect 430 171 437 173
rect 443 182 450 184
rect 443 180 445 182
rect 447 180 450 182
rect 443 175 450 180
rect 443 173 445 175
rect 447 173 450 175
rect 443 171 450 173
rect 430 156 435 171
rect 445 156 450 171
rect 452 167 460 184
rect 452 165 455 167
rect 457 165 460 167
rect 452 160 460 165
rect 452 158 455 160
rect 457 158 460 160
rect 452 156 460 158
rect 462 175 470 184
rect 462 173 465 175
rect 467 173 470 175
rect 462 168 470 173
rect 462 166 465 168
rect 467 166 470 168
rect 462 156 470 166
rect 472 167 488 184
rect 472 165 477 167
rect 479 165 488 167
rect 472 160 488 165
rect 472 158 477 160
rect 479 159 488 160
rect 490 159 495 184
rect 497 181 502 184
rect 497 179 505 181
rect 497 177 500 179
rect 502 177 505 179
rect 497 168 505 177
rect 507 168 518 181
rect 497 159 502 168
rect 509 160 518 168
rect 479 158 486 159
rect 472 156 486 158
rect 509 158 512 160
rect 514 158 518 160
rect 509 156 518 158
rect 520 179 527 181
rect 520 177 523 179
rect 525 177 527 179
rect 551 177 559 184
rect 520 172 527 177
rect 520 170 523 172
rect 525 170 527 172
rect 520 168 527 170
rect 534 169 539 177
rect 520 156 525 168
rect 532 167 539 169
rect 532 165 534 167
rect 536 165 539 167
rect 532 163 539 165
rect 534 156 539 163
rect 541 156 546 177
rect 548 166 559 177
rect 561 179 566 184
rect 561 177 568 179
rect 561 175 564 177
rect 566 175 568 177
rect 601 176 607 183
rect 561 170 568 175
rect 561 168 564 170
rect 566 168 568 170
rect 561 166 568 168
rect 580 167 587 176
rect 548 160 557 166
rect 580 165 582 167
rect 584 165 587 167
rect 580 163 587 165
rect 589 174 597 176
rect 589 172 592 174
rect 594 172 597 174
rect 589 167 597 172
rect 589 165 592 167
rect 594 165 597 167
rect 589 163 597 165
rect 599 169 607 176
rect 599 167 602 169
rect 604 167 607 169
rect 599 165 607 167
rect 609 181 616 183
rect 645 181 650 184
rect 609 179 612 181
rect 614 179 616 181
rect 609 174 616 179
rect 609 172 612 174
rect 614 172 616 174
rect 609 170 616 172
rect 620 179 627 181
rect 620 177 622 179
rect 624 177 627 179
rect 620 172 627 177
rect 620 170 622 172
rect 624 170 627 172
rect 609 165 614 170
rect 620 168 627 170
rect 599 163 605 165
rect 548 158 553 160
rect 555 158 557 160
rect 548 156 557 158
rect 622 156 627 168
rect 629 168 640 181
rect 642 179 650 181
rect 642 177 645 179
rect 647 177 650 179
rect 642 168 650 177
rect 629 160 638 168
rect 629 158 633 160
rect 635 158 638 160
rect 645 159 650 168
rect 652 159 657 184
rect 659 167 675 184
rect 659 165 668 167
rect 670 165 675 167
rect 659 160 675 165
rect 659 159 668 160
rect 629 156 638 158
rect 661 158 668 159
rect 670 158 675 160
rect 661 156 675 158
rect 677 175 685 184
rect 677 173 680 175
rect 682 173 685 175
rect 677 168 685 173
rect 677 166 680 168
rect 682 166 685 168
rect 677 156 685 166
rect 687 167 695 184
rect 687 165 690 167
rect 692 165 695 167
rect 687 160 695 165
rect 687 158 690 160
rect 692 158 695 160
rect 687 156 695 158
rect 697 182 704 184
rect 697 180 700 182
rect 702 180 704 182
rect 697 175 704 180
rect 697 173 700 175
rect 702 173 704 175
rect 697 171 704 173
rect 710 182 717 184
rect 710 180 712 182
rect 714 180 717 182
rect 710 175 717 180
rect 710 173 712 175
rect 714 173 717 175
rect 710 171 717 173
rect 697 156 702 171
rect 712 156 717 171
rect 719 167 727 184
rect 719 165 722 167
rect 724 165 727 167
rect 719 160 727 165
rect 719 158 722 160
rect 724 158 727 160
rect 719 156 727 158
rect 729 175 737 184
rect 729 173 732 175
rect 734 173 737 175
rect 729 168 737 173
rect 729 166 732 168
rect 734 166 737 168
rect 729 156 737 166
rect 739 167 755 184
rect 739 165 744 167
rect 746 165 755 167
rect 739 160 755 165
rect 739 158 744 160
rect 746 159 755 160
rect 757 159 762 184
rect 764 181 769 184
rect 764 179 772 181
rect 764 177 767 179
rect 769 177 772 179
rect 764 168 772 177
rect 774 168 785 181
rect 764 159 769 168
rect 776 160 785 168
rect 746 158 753 159
rect 739 156 753 158
rect 776 158 779 160
rect 781 158 785 160
rect 776 156 785 158
rect 787 179 794 181
rect 787 177 790 179
rect 792 177 794 179
rect 818 177 826 184
rect 787 172 794 177
rect 787 170 790 172
rect 792 170 794 172
rect 787 168 794 170
rect 801 169 806 177
rect 787 156 792 168
rect 799 167 806 169
rect 799 165 801 167
rect 803 165 806 167
rect 799 163 806 165
rect 801 156 806 163
rect 808 156 813 177
rect 815 166 826 177
rect 828 179 833 184
rect 828 177 835 179
rect 828 175 831 177
rect 833 175 835 177
rect 828 170 835 175
rect 828 168 831 170
rect 833 168 835 170
rect 828 166 835 168
rect 815 160 824 166
rect 815 158 820 160
rect 822 158 824 160
rect 815 156 824 158
rect 6 135 13 137
rect 6 133 8 135
rect 10 133 13 135
rect 6 124 13 133
rect 15 135 23 137
rect 15 133 18 135
rect 20 133 23 135
rect 15 128 23 133
rect 15 126 18 128
rect 20 126 23 128
rect 15 124 23 126
rect 25 135 31 137
rect 46 135 53 137
rect 25 133 33 135
rect 25 131 28 133
rect 30 131 33 133
rect 25 124 33 131
rect 27 117 33 124
rect 35 133 40 135
rect 46 133 48 135
rect 50 133 53 135
rect 35 131 42 133
rect 35 129 38 131
rect 40 129 42 131
rect 35 123 42 129
rect 46 124 53 133
rect 55 135 63 137
rect 55 133 58 135
rect 60 133 63 135
rect 55 128 63 133
rect 55 126 58 128
rect 60 126 63 128
rect 55 124 63 126
rect 65 135 71 137
rect 65 133 73 135
rect 65 131 68 133
rect 70 131 73 133
rect 65 124 73 131
rect 35 121 38 123
rect 40 121 42 123
rect 35 117 42 121
rect 67 117 73 124
rect 75 130 80 135
rect 88 132 93 144
rect 86 130 93 132
rect 75 128 82 130
rect 75 126 78 128
rect 80 126 82 128
rect 75 121 82 126
rect 75 119 78 121
rect 80 119 82 121
rect 86 128 88 130
rect 90 128 93 130
rect 86 123 93 128
rect 86 121 88 123
rect 90 121 93 123
rect 86 119 93 121
rect 95 142 104 144
rect 95 140 99 142
rect 101 140 104 142
rect 127 142 141 144
rect 127 141 134 142
rect 95 132 104 140
rect 111 132 116 141
rect 95 119 106 132
rect 108 123 116 132
rect 108 121 111 123
rect 113 121 116 123
rect 108 119 116 121
rect 75 117 82 119
rect 111 116 116 119
rect 118 116 123 141
rect 125 140 134 141
rect 136 140 141 142
rect 125 135 141 140
rect 125 133 134 135
rect 136 133 141 135
rect 125 116 141 133
rect 143 134 151 144
rect 143 132 146 134
rect 148 132 151 134
rect 143 127 151 132
rect 143 125 146 127
rect 148 125 151 127
rect 143 116 151 125
rect 153 142 161 144
rect 153 140 156 142
rect 158 140 161 142
rect 153 135 161 140
rect 153 133 156 135
rect 158 133 161 135
rect 153 116 161 133
rect 163 129 168 144
rect 178 129 183 144
rect 163 127 170 129
rect 163 125 166 127
rect 168 125 170 127
rect 163 120 170 125
rect 163 118 166 120
rect 168 118 170 120
rect 163 116 170 118
rect 176 127 183 129
rect 176 125 178 127
rect 180 125 183 127
rect 176 120 183 125
rect 176 118 178 120
rect 180 118 183 120
rect 176 116 183 118
rect 185 142 193 144
rect 185 140 188 142
rect 190 140 193 142
rect 185 135 193 140
rect 185 133 188 135
rect 190 133 193 135
rect 185 116 193 133
rect 195 134 203 144
rect 195 132 198 134
rect 200 132 203 134
rect 195 127 203 132
rect 195 125 198 127
rect 200 125 203 127
rect 195 116 203 125
rect 205 142 219 144
rect 205 140 210 142
rect 212 141 219 142
rect 242 142 251 144
rect 212 140 221 141
rect 205 135 221 140
rect 205 133 210 135
rect 212 133 221 135
rect 205 116 221 133
rect 223 116 228 141
rect 230 132 235 141
rect 242 140 245 142
rect 247 140 251 142
rect 242 132 251 140
rect 230 123 238 132
rect 230 121 233 123
rect 235 121 238 123
rect 230 119 238 121
rect 240 119 251 132
rect 253 132 258 144
rect 267 137 272 144
rect 265 135 272 137
rect 265 133 267 135
rect 269 133 272 135
rect 253 130 260 132
rect 265 131 272 133
rect 253 128 256 130
rect 258 128 260 130
rect 253 123 260 128
rect 267 123 272 131
rect 274 123 279 144
rect 281 142 290 144
rect 281 140 286 142
rect 288 140 290 142
rect 281 134 290 140
rect 313 135 320 137
rect 281 123 292 134
rect 253 121 256 123
rect 258 121 260 123
rect 253 119 260 121
rect 230 116 235 119
rect 284 116 292 123
rect 294 132 301 134
rect 294 130 297 132
rect 299 130 301 132
rect 294 125 301 130
rect 294 123 297 125
rect 299 123 301 125
rect 313 133 315 135
rect 317 133 320 135
rect 313 124 320 133
rect 322 135 330 137
rect 322 133 325 135
rect 327 133 330 135
rect 322 128 330 133
rect 322 126 325 128
rect 327 126 330 128
rect 322 124 330 126
rect 332 135 338 137
rect 332 133 340 135
rect 332 131 335 133
rect 337 131 340 133
rect 332 124 340 131
rect 294 121 301 123
rect 294 116 299 121
rect 334 117 340 124
rect 342 130 347 135
rect 355 132 360 144
rect 353 130 360 132
rect 342 128 349 130
rect 342 126 345 128
rect 347 126 349 128
rect 342 121 349 126
rect 342 119 345 121
rect 347 119 349 121
rect 353 128 355 130
rect 357 128 360 130
rect 353 123 360 128
rect 353 121 355 123
rect 357 121 360 123
rect 353 119 360 121
rect 362 142 371 144
rect 362 140 366 142
rect 368 140 371 142
rect 394 142 408 144
rect 394 141 401 142
rect 362 132 371 140
rect 378 132 383 141
rect 362 119 373 132
rect 375 123 383 132
rect 375 121 378 123
rect 380 121 383 123
rect 375 119 383 121
rect 342 117 349 119
rect 378 116 383 119
rect 385 116 390 141
rect 392 140 401 141
rect 403 140 408 142
rect 392 135 408 140
rect 392 133 401 135
rect 403 133 408 135
rect 392 116 408 133
rect 410 134 418 144
rect 410 132 413 134
rect 415 132 418 134
rect 410 127 418 132
rect 410 125 413 127
rect 415 125 418 127
rect 410 116 418 125
rect 420 142 428 144
rect 420 140 423 142
rect 425 140 428 142
rect 420 135 428 140
rect 420 133 423 135
rect 425 133 428 135
rect 420 116 428 133
rect 430 129 435 144
rect 445 129 450 144
rect 430 127 437 129
rect 430 125 433 127
rect 435 125 437 127
rect 430 120 437 125
rect 430 118 433 120
rect 435 118 437 120
rect 430 116 437 118
rect 443 127 450 129
rect 443 125 445 127
rect 447 125 450 127
rect 443 120 450 125
rect 443 118 445 120
rect 447 118 450 120
rect 443 116 450 118
rect 452 142 460 144
rect 452 140 455 142
rect 457 140 460 142
rect 452 135 460 140
rect 452 133 455 135
rect 457 133 460 135
rect 452 116 460 133
rect 462 134 470 144
rect 462 132 465 134
rect 467 132 470 134
rect 462 127 470 132
rect 462 125 465 127
rect 467 125 470 127
rect 462 116 470 125
rect 472 142 486 144
rect 472 140 477 142
rect 479 141 486 142
rect 509 142 518 144
rect 479 140 488 141
rect 472 135 488 140
rect 472 133 477 135
rect 479 133 488 135
rect 472 116 488 133
rect 490 116 495 141
rect 497 132 502 141
rect 509 140 512 142
rect 514 140 518 142
rect 509 132 518 140
rect 497 123 505 132
rect 497 121 500 123
rect 502 121 505 123
rect 497 119 505 121
rect 507 119 518 132
rect 520 132 525 144
rect 534 137 539 144
rect 532 135 539 137
rect 532 133 534 135
rect 536 133 539 135
rect 520 130 527 132
rect 532 131 539 133
rect 520 128 523 130
rect 525 128 527 130
rect 520 123 527 128
rect 534 123 539 131
rect 541 123 546 144
rect 548 142 557 144
rect 548 140 553 142
rect 555 140 557 142
rect 548 134 557 140
rect 580 135 587 137
rect 548 123 559 134
rect 520 121 523 123
rect 525 121 527 123
rect 520 119 527 121
rect 497 116 502 119
rect 551 116 559 123
rect 561 132 568 134
rect 561 130 564 132
rect 566 130 568 132
rect 561 125 568 130
rect 561 123 564 125
rect 566 123 568 125
rect 580 133 582 135
rect 584 133 587 135
rect 580 124 587 133
rect 589 135 597 137
rect 589 133 592 135
rect 594 133 597 135
rect 589 128 597 133
rect 589 126 592 128
rect 594 126 597 128
rect 589 124 597 126
rect 599 135 605 137
rect 599 133 607 135
rect 599 131 602 133
rect 604 131 607 133
rect 599 124 607 131
rect 561 121 568 123
rect 561 116 566 121
rect 601 117 607 124
rect 609 130 614 135
rect 622 132 627 144
rect 620 130 627 132
rect 609 128 616 130
rect 609 126 612 128
rect 614 126 616 128
rect 609 121 616 126
rect 609 119 612 121
rect 614 119 616 121
rect 620 128 622 130
rect 624 128 627 130
rect 620 123 627 128
rect 620 121 622 123
rect 624 121 627 123
rect 620 119 627 121
rect 629 142 638 144
rect 629 140 633 142
rect 635 140 638 142
rect 661 142 675 144
rect 661 141 668 142
rect 629 132 638 140
rect 645 132 650 141
rect 629 119 640 132
rect 642 123 650 132
rect 642 121 645 123
rect 647 121 650 123
rect 642 119 650 121
rect 609 117 616 119
rect 645 116 650 119
rect 652 116 657 141
rect 659 140 668 141
rect 670 140 675 142
rect 659 135 675 140
rect 659 133 668 135
rect 670 133 675 135
rect 659 116 675 133
rect 677 134 685 144
rect 677 132 680 134
rect 682 132 685 134
rect 677 127 685 132
rect 677 125 680 127
rect 682 125 685 127
rect 677 116 685 125
rect 687 142 695 144
rect 687 140 690 142
rect 692 140 695 142
rect 687 135 695 140
rect 687 133 690 135
rect 692 133 695 135
rect 687 116 695 133
rect 697 129 702 144
rect 712 129 717 144
rect 697 127 704 129
rect 697 125 700 127
rect 702 125 704 127
rect 697 120 704 125
rect 697 118 700 120
rect 702 118 704 120
rect 697 116 704 118
rect 710 127 717 129
rect 710 125 712 127
rect 714 125 717 127
rect 710 120 717 125
rect 710 118 712 120
rect 714 118 717 120
rect 710 116 717 118
rect 719 142 727 144
rect 719 140 722 142
rect 724 140 727 142
rect 719 135 727 140
rect 719 133 722 135
rect 724 133 727 135
rect 719 116 727 133
rect 729 134 737 144
rect 729 132 732 134
rect 734 132 737 134
rect 729 127 737 132
rect 729 125 732 127
rect 734 125 737 127
rect 729 116 737 125
rect 739 142 753 144
rect 739 140 744 142
rect 746 141 753 142
rect 776 142 785 144
rect 746 140 755 141
rect 739 135 755 140
rect 739 133 744 135
rect 746 133 755 135
rect 739 116 755 133
rect 757 116 762 141
rect 764 132 769 141
rect 776 140 779 142
rect 781 140 785 142
rect 776 132 785 140
rect 764 123 772 132
rect 764 121 767 123
rect 769 121 772 123
rect 764 119 772 121
rect 774 119 785 132
rect 787 132 792 144
rect 801 137 806 144
rect 799 135 806 137
rect 799 133 801 135
rect 803 133 806 135
rect 787 130 794 132
rect 799 131 806 133
rect 787 128 790 130
rect 792 128 794 130
rect 787 123 794 128
rect 801 123 806 131
rect 808 123 813 144
rect 815 142 824 144
rect 815 140 820 142
rect 822 140 824 142
rect 815 134 824 140
rect 815 123 826 134
rect 787 121 790 123
rect 792 121 794 123
rect 787 119 794 121
rect 764 116 769 119
rect 818 116 826 123
rect 828 132 835 134
rect 828 130 831 132
rect 833 130 835 132
rect 828 125 835 130
rect 828 123 831 125
rect 833 123 835 125
rect 828 121 835 123
rect 828 116 833 121
rect 27 32 33 39
rect 6 23 13 32
rect 6 21 8 23
rect 10 21 13 23
rect 6 19 13 21
rect 15 30 23 32
rect 15 28 18 30
rect 20 28 23 30
rect 15 23 23 28
rect 15 21 18 23
rect 20 21 23 23
rect 15 19 23 21
rect 25 25 33 32
rect 25 23 28 25
rect 30 23 33 25
rect 25 21 33 23
rect 35 37 42 39
rect 35 35 38 37
rect 40 35 42 37
rect 35 30 42 35
rect 67 32 73 39
rect 35 28 38 30
rect 40 28 42 30
rect 35 26 42 28
rect 35 21 40 26
rect 46 23 53 32
rect 46 21 48 23
rect 50 21 53 23
rect 25 19 31 21
rect 46 19 53 21
rect 55 30 63 32
rect 55 28 58 30
rect 60 28 63 30
rect 55 23 63 28
rect 55 21 58 23
rect 60 21 63 23
rect 55 19 63 21
rect 65 25 73 32
rect 65 23 68 25
rect 70 23 73 25
rect 65 21 73 23
rect 75 37 82 39
rect 111 37 116 40
rect 75 35 78 37
rect 80 35 82 37
rect 75 30 82 35
rect 75 28 78 30
rect 80 28 82 30
rect 75 26 82 28
rect 86 35 93 37
rect 86 33 88 35
rect 90 33 93 35
rect 86 28 93 33
rect 86 26 88 28
rect 90 26 93 28
rect 75 21 80 26
rect 86 24 93 26
rect 65 19 71 21
rect 88 12 93 24
rect 95 24 106 37
rect 108 35 116 37
rect 108 33 111 35
rect 113 33 116 35
rect 108 24 116 33
rect 95 16 104 24
rect 95 14 99 16
rect 101 14 104 16
rect 111 15 116 24
rect 118 15 123 40
rect 125 23 141 40
rect 125 21 134 23
rect 136 21 141 23
rect 125 16 141 21
rect 125 15 134 16
rect 95 12 104 14
rect 127 14 134 15
rect 136 14 141 16
rect 127 12 141 14
rect 143 31 151 40
rect 143 29 146 31
rect 148 29 151 31
rect 143 24 151 29
rect 143 22 146 24
rect 148 22 151 24
rect 143 12 151 22
rect 153 23 161 40
rect 153 21 156 23
rect 158 21 161 23
rect 153 16 161 21
rect 153 14 156 16
rect 158 14 161 16
rect 153 12 161 14
rect 163 38 170 40
rect 163 36 166 38
rect 168 36 170 38
rect 163 31 170 36
rect 163 29 166 31
rect 168 29 170 31
rect 163 27 170 29
rect 176 38 183 40
rect 176 36 178 38
rect 180 36 183 38
rect 176 31 183 36
rect 176 29 178 31
rect 180 29 183 31
rect 176 27 183 29
rect 163 12 168 27
rect 178 12 183 27
rect 185 23 193 40
rect 185 21 188 23
rect 190 21 193 23
rect 185 16 193 21
rect 185 14 188 16
rect 190 14 193 16
rect 185 12 193 14
rect 195 31 203 40
rect 195 29 198 31
rect 200 29 203 31
rect 195 24 203 29
rect 195 22 198 24
rect 200 22 203 24
rect 195 12 203 22
rect 205 23 221 40
rect 205 21 210 23
rect 212 21 221 23
rect 205 16 221 21
rect 205 14 210 16
rect 212 15 221 16
rect 223 15 228 40
rect 230 37 235 40
rect 230 35 238 37
rect 230 33 233 35
rect 235 33 238 35
rect 230 24 238 33
rect 240 24 251 37
rect 230 15 235 24
rect 242 16 251 24
rect 212 14 219 15
rect 205 12 219 14
rect 242 14 245 16
rect 247 14 251 16
rect 242 12 251 14
rect 253 35 260 37
rect 253 33 256 35
rect 258 33 260 35
rect 284 33 292 40
rect 253 28 260 33
rect 253 26 256 28
rect 258 26 260 28
rect 253 24 260 26
rect 267 25 272 33
rect 253 12 258 24
rect 265 23 272 25
rect 265 21 267 23
rect 269 21 272 23
rect 265 19 272 21
rect 267 12 272 19
rect 274 12 279 33
rect 281 22 292 33
rect 294 35 299 40
rect 294 33 301 35
rect 294 31 297 33
rect 299 31 301 33
rect 334 32 340 39
rect 294 26 301 31
rect 294 24 297 26
rect 299 24 301 26
rect 294 22 301 24
rect 313 23 320 32
rect 281 16 290 22
rect 313 21 315 23
rect 317 21 320 23
rect 313 19 320 21
rect 322 30 330 32
rect 322 28 325 30
rect 327 28 330 30
rect 322 23 330 28
rect 322 21 325 23
rect 327 21 330 23
rect 322 19 330 21
rect 332 25 340 32
rect 332 23 335 25
rect 337 23 340 25
rect 332 21 340 23
rect 342 37 349 39
rect 378 37 383 40
rect 342 35 345 37
rect 347 35 349 37
rect 342 30 349 35
rect 342 28 345 30
rect 347 28 349 30
rect 342 26 349 28
rect 353 35 360 37
rect 353 33 355 35
rect 357 33 360 35
rect 353 28 360 33
rect 353 26 355 28
rect 357 26 360 28
rect 342 21 347 26
rect 353 24 360 26
rect 332 19 338 21
rect 281 14 286 16
rect 288 14 290 16
rect 281 12 290 14
rect 355 12 360 24
rect 362 24 373 37
rect 375 35 383 37
rect 375 33 378 35
rect 380 33 383 35
rect 375 24 383 33
rect 362 16 371 24
rect 362 14 366 16
rect 368 14 371 16
rect 378 15 383 24
rect 385 15 390 40
rect 392 23 408 40
rect 392 21 401 23
rect 403 21 408 23
rect 392 16 408 21
rect 392 15 401 16
rect 362 12 371 14
rect 394 14 401 15
rect 403 14 408 16
rect 394 12 408 14
rect 410 31 418 40
rect 410 29 413 31
rect 415 29 418 31
rect 410 24 418 29
rect 410 22 413 24
rect 415 22 418 24
rect 410 12 418 22
rect 420 23 428 40
rect 420 21 423 23
rect 425 21 428 23
rect 420 16 428 21
rect 420 14 423 16
rect 425 14 428 16
rect 420 12 428 14
rect 430 38 437 40
rect 430 36 433 38
rect 435 36 437 38
rect 430 31 437 36
rect 430 29 433 31
rect 435 29 437 31
rect 430 27 437 29
rect 443 38 450 40
rect 443 36 445 38
rect 447 36 450 38
rect 443 31 450 36
rect 443 29 445 31
rect 447 29 450 31
rect 443 27 450 29
rect 430 12 435 27
rect 445 12 450 27
rect 452 23 460 40
rect 452 21 455 23
rect 457 21 460 23
rect 452 16 460 21
rect 452 14 455 16
rect 457 14 460 16
rect 452 12 460 14
rect 462 31 470 40
rect 462 29 465 31
rect 467 29 470 31
rect 462 24 470 29
rect 462 22 465 24
rect 467 22 470 24
rect 462 12 470 22
rect 472 23 488 40
rect 472 21 477 23
rect 479 21 488 23
rect 472 16 488 21
rect 472 14 477 16
rect 479 15 488 16
rect 490 15 495 40
rect 497 37 502 40
rect 497 35 505 37
rect 497 33 500 35
rect 502 33 505 35
rect 497 24 505 33
rect 507 24 518 37
rect 497 15 502 24
rect 509 16 518 24
rect 479 14 486 15
rect 472 12 486 14
rect 509 14 512 16
rect 514 14 518 16
rect 509 12 518 14
rect 520 35 527 37
rect 520 33 523 35
rect 525 33 527 35
rect 551 33 559 40
rect 520 28 527 33
rect 520 26 523 28
rect 525 26 527 28
rect 520 24 527 26
rect 534 25 539 33
rect 520 12 525 24
rect 532 23 539 25
rect 532 21 534 23
rect 536 21 539 23
rect 532 19 539 21
rect 534 12 539 19
rect 541 12 546 33
rect 548 22 559 33
rect 561 35 566 40
rect 561 33 568 35
rect 561 31 564 33
rect 566 31 568 33
rect 601 32 607 39
rect 561 26 568 31
rect 561 24 564 26
rect 566 24 568 26
rect 561 22 568 24
rect 580 23 587 32
rect 548 16 557 22
rect 580 21 582 23
rect 584 21 587 23
rect 580 19 587 21
rect 589 30 597 32
rect 589 28 592 30
rect 594 28 597 30
rect 589 23 597 28
rect 589 21 592 23
rect 594 21 597 23
rect 589 19 597 21
rect 599 25 607 32
rect 599 23 602 25
rect 604 23 607 25
rect 599 21 607 23
rect 609 37 616 39
rect 645 37 650 40
rect 609 35 612 37
rect 614 35 616 37
rect 609 30 616 35
rect 609 28 612 30
rect 614 28 616 30
rect 609 26 616 28
rect 620 35 627 37
rect 620 33 622 35
rect 624 33 627 35
rect 620 28 627 33
rect 620 26 622 28
rect 624 26 627 28
rect 609 21 614 26
rect 620 24 627 26
rect 599 19 605 21
rect 548 14 553 16
rect 555 14 557 16
rect 548 12 557 14
rect 622 12 627 24
rect 629 24 640 37
rect 642 35 650 37
rect 642 33 645 35
rect 647 33 650 35
rect 642 24 650 33
rect 629 16 638 24
rect 629 14 633 16
rect 635 14 638 16
rect 645 15 650 24
rect 652 15 657 40
rect 659 23 675 40
rect 659 21 668 23
rect 670 21 675 23
rect 659 16 675 21
rect 659 15 668 16
rect 629 12 638 14
rect 661 14 668 15
rect 670 14 675 16
rect 661 12 675 14
rect 677 31 685 40
rect 677 29 680 31
rect 682 29 685 31
rect 677 24 685 29
rect 677 22 680 24
rect 682 22 685 24
rect 677 12 685 22
rect 687 23 695 40
rect 687 21 690 23
rect 692 21 695 23
rect 687 16 695 21
rect 687 14 690 16
rect 692 14 695 16
rect 687 12 695 14
rect 697 38 704 40
rect 697 36 700 38
rect 702 36 704 38
rect 697 31 704 36
rect 697 29 700 31
rect 702 29 704 31
rect 697 27 704 29
rect 710 38 717 40
rect 710 36 712 38
rect 714 36 717 38
rect 710 31 717 36
rect 710 29 712 31
rect 714 29 717 31
rect 710 27 717 29
rect 697 12 702 27
rect 712 12 717 27
rect 719 23 727 40
rect 719 21 722 23
rect 724 21 727 23
rect 719 16 727 21
rect 719 14 722 16
rect 724 14 727 16
rect 719 12 727 14
rect 729 31 737 40
rect 729 29 732 31
rect 734 29 737 31
rect 729 24 737 29
rect 729 22 732 24
rect 734 22 737 24
rect 729 12 737 22
rect 739 23 755 40
rect 739 21 744 23
rect 746 21 755 23
rect 739 16 755 21
rect 739 14 744 16
rect 746 15 755 16
rect 757 15 762 40
rect 764 37 769 40
rect 764 35 772 37
rect 764 33 767 35
rect 769 33 772 35
rect 764 24 772 33
rect 774 24 785 37
rect 764 15 769 24
rect 776 16 785 24
rect 746 14 753 15
rect 739 12 753 14
rect 776 14 779 16
rect 781 14 785 16
rect 776 12 785 14
rect 787 35 794 37
rect 787 33 790 35
rect 792 33 794 35
rect 818 33 826 40
rect 787 28 794 33
rect 787 26 790 28
rect 792 26 794 28
rect 787 24 794 26
rect 801 25 806 33
rect 787 12 792 24
rect 799 23 806 25
rect 799 21 801 23
rect 803 21 806 23
rect 799 19 806 21
rect 801 12 806 19
rect 808 12 813 33
rect 815 22 826 33
rect 828 35 833 40
rect 828 33 835 35
rect 828 31 831 33
rect 833 31 835 33
rect 828 26 835 31
rect 828 24 831 26
rect 833 24 835 26
rect 828 22 835 24
rect 815 16 824 22
rect 815 14 820 16
rect 822 14 824 16
rect 815 12 824 14
rect 434 -21 439 0
rect 432 -23 439 -21
rect 432 -25 434 -23
rect 436 -25 439 -23
rect 432 -27 439 -25
rect 441 -2 453 0
rect 441 -4 444 -2
rect 446 -4 453 -2
rect 441 -9 453 -4
rect 470 -9 475 0
rect 441 -11 444 -9
rect 446 -11 455 -9
rect 441 -27 455 -11
rect 457 -16 465 -9
rect 457 -18 460 -16
rect 462 -18 465 -16
rect 457 -23 465 -18
rect 457 -25 460 -23
rect 462 -25 465 -23
rect 457 -27 465 -25
rect 467 -16 475 -9
rect 467 -18 470 -16
rect 472 -18 475 -16
rect 467 -27 475 -18
rect 477 -6 482 0
rect 477 -8 484 -6
rect 477 -10 480 -8
rect 482 -10 484 -8
rect 477 -12 484 -10
rect 490 -12 495 0
rect 477 -27 482 -12
rect 488 -14 495 -12
rect 488 -16 490 -14
rect 492 -16 495 -14
rect 488 -21 495 -16
rect 488 -23 490 -21
rect 492 -23 495 -21
rect 488 -25 495 -23
rect 497 -2 506 0
rect 497 -4 501 -2
rect 503 -4 506 -2
rect 529 -2 543 0
rect 529 -3 536 -2
rect 497 -12 506 -4
rect 513 -12 518 -3
rect 497 -25 508 -12
rect 510 -21 518 -12
rect 510 -23 513 -21
rect 515 -23 518 -21
rect 510 -25 518 -23
rect 513 -28 518 -25
rect 520 -28 525 -3
rect 527 -4 536 -3
rect 538 -4 543 -2
rect 527 -9 543 -4
rect 527 -11 536 -9
rect 538 -11 543 -9
rect 527 -28 543 -11
rect 545 -10 553 0
rect 545 -12 548 -10
rect 550 -12 553 -10
rect 545 -17 553 -12
rect 545 -19 548 -17
rect 550 -19 553 -17
rect 545 -28 553 -19
rect 555 -2 563 0
rect 555 -4 558 -2
rect 560 -4 563 -2
rect 555 -9 563 -4
rect 555 -11 558 -9
rect 560 -11 563 -9
rect 555 -28 563 -11
rect 565 -15 570 0
rect 580 -15 585 0
rect 565 -17 572 -15
rect 565 -19 568 -17
rect 570 -19 572 -17
rect 565 -24 572 -19
rect 565 -26 568 -24
rect 570 -26 572 -24
rect 565 -28 572 -26
rect 578 -17 585 -15
rect 578 -19 580 -17
rect 582 -19 585 -17
rect 578 -24 585 -19
rect 578 -26 580 -24
rect 582 -26 585 -24
rect 578 -28 585 -26
rect 587 -2 595 0
rect 587 -4 590 -2
rect 592 -4 595 -2
rect 587 -9 595 -4
rect 587 -11 590 -9
rect 592 -11 595 -9
rect 587 -28 595 -11
rect 597 -10 605 0
rect 597 -12 600 -10
rect 602 -12 605 -10
rect 597 -17 605 -12
rect 597 -19 600 -17
rect 602 -19 605 -17
rect 597 -28 605 -19
rect 607 -2 621 0
rect 607 -4 612 -2
rect 614 -3 621 -2
rect 644 -2 653 0
rect 614 -4 623 -3
rect 607 -9 623 -4
rect 607 -11 612 -9
rect 614 -11 623 -9
rect 607 -28 623 -11
rect 625 -28 630 -3
rect 632 -12 637 -3
rect 644 -4 647 -2
rect 649 -4 653 -2
rect 644 -12 653 -4
rect 632 -21 640 -12
rect 632 -23 635 -21
rect 637 -23 640 -21
rect 632 -25 640 -23
rect 642 -25 653 -12
rect 655 -12 660 0
rect 669 -7 674 0
rect 667 -9 674 -7
rect 667 -11 669 -9
rect 671 -11 674 -9
rect 655 -14 662 -12
rect 667 -13 674 -11
rect 655 -16 658 -14
rect 660 -16 662 -14
rect 655 -21 662 -16
rect 669 -21 674 -13
rect 676 -21 681 0
rect 683 -2 692 0
rect 683 -4 688 -2
rect 690 -4 692 -2
rect 720 -2 727 0
rect 683 -10 692 -4
rect 720 -4 722 -2
rect 724 -4 727 -2
rect 683 -21 694 -10
rect 655 -23 658 -21
rect 660 -23 662 -21
rect 655 -25 662 -23
rect 632 -28 637 -25
rect 686 -28 694 -21
rect 696 -12 703 -10
rect 696 -14 699 -12
rect 701 -14 703 -12
rect 696 -19 703 -14
rect 720 -12 727 -4
rect 696 -21 699 -19
rect 701 -21 703 -19
rect 721 -16 727 -12
rect 729 -16 734 0
rect 736 -12 744 0
rect 736 -14 739 -12
rect 741 -14 744 -12
rect 736 -16 744 -14
rect 746 -16 751 0
rect 753 -2 761 0
rect 753 -4 756 -2
rect 758 -4 761 -2
rect 753 -16 761 -4
rect 721 -20 725 -16
rect 696 -23 703 -21
rect 712 -22 717 -20
rect 696 -28 701 -23
rect 710 -24 717 -22
rect 710 -26 712 -24
rect 714 -26 717 -24
rect 710 -28 717 -26
rect 719 -28 725 -20
rect 756 -18 761 -16
rect 763 -7 768 0
rect 784 -2 791 0
rect 784 -4 786 -2
rect 788 -4 791 -2
rect 763 -9 770 -7
rect 763 -11 766 -9
rect 768 -11 770 -9
rect 763 -13 770 -11
rect 784 -12 791 -4
rect 763 -18 768 -13
rect 785 -16 791 -12
rect 793 -16 798 0
rect 800 -12 808 0
rect 800 -14 803 -12
rect 805 -14 808 -12
rect 800 -16 808 -14
rect 810 -16 815 0
rect 817 -2 825 0
rect 817 -4 820 -2
rect 822 -4 825 -2
rect 817 -16 825 -4
rect 785 -20 789 -16
rect 776 -22 781 -20
rect 774 -24 781 -22
rect 774 -26 776 -24
rect 778 -26 781 -24
rect 774 -28 781 -26
rect 783 -28 789 -20
rect 820 -18 825 -16
rect 827 -7 832 0
rect 827 -9 834 -7
rect 827 -11 830 -9
rect 832 -11 834 -9
rect 827 -13 834 -11
rect 827 -18 832 -13
rect 432 -107 439 -105
rect 432 -109 434 -107
rect 436 -109 439 -107
rect 432 -111 439 -109
rect 434 -132 439 -111
rect 441 -121 455 -105
rect 441 -123 444 -121
rect 446 -123 455 -121
rect 457 -107 465 -105
rect 457 -109 460 -107
rect 462 -109 465 -107
rect 457 -114 465 -109
rect 457 -116 460 -114
rect 462 -116 465 -114
rect 457 -123 465 -116
rect 467 -114 475 -105
rect 467 -116 470 -114
rect 472 -116 475 -114
rect 467 -123 475 -116
rect 441 -128 453 -123
rect 441 -130 444 -128
rect 446 -130 453 -128
rect 441 -132 453 -130
rect 470 -132 475 -123
rect 477 -120 482 -105
rect 513 -107 518 -104
rect 488 -109 495 -107
rect 488 -111 490 -109
rect 492 -111 495 -109
rect 488 -116 495 -111
rect 488 -118 490 -116
rect 492 -118 495 -116
rect 488 -120 495 -118
rect 477 -122 484 -120
rect 477 -124 480 -122
rect 482 -124 484 -122
rect 477 -126 484 -124
rect 477 -132 482 -126
rect 490 -132 495 -120
rect 497 -120 508 -107
rect 510 -109 518 -107
rect 510 -111 513 -109
rect 515 -111 518 -109
rect 510 -120 518 -111
rect 497 -128 506 -120
rect 497 -130 501 -128
rect 503 -130 506 -128
rect 513 -129 518 -120
rect 520 -129 525 -104
rect 527 -121 543 -104
rect 527 -123 536 -121
rect 538 -123 543 -121
rect 527 -128 543 -123
rect 527 -129 536 -128
rect 497 -132 506 -130
rect 529 -130 536 -129
rect 538 -130 543 -128
rect 529 -132 543 -130
rect 545 -113 553 -104
rect 545 -115 548 -113
rect 550 -115 553 -113
rect 545 -120 553 -115
rect 545 -122 548 -120
rect 550 -122 553 -120
rect 545 -132 553 -122
rect 555 -121 563 -104
rect 555 -123 558 -121
rect 560 -123 563 -121
rect 555 -128 563 -123
rect 555 -130 558 -128
rect 560 -130 563 -128
rect 555 -132 563 -130
rect 565 -106 572 -104
rect 565 -108 568 -106
rect 570 -108 572 -106
rect 565 -113 572 -108
rect 565 -115 568 -113
rect 570 -115 572 -113
rect 565 -117 572 -115
rect 578 -106 585 -104
rect 578 -108 580 -106
rect 582 -108 585 -106
rect 578 -113 585 -108
rect 578 -115 580 -113
rect 582 -115 585 -113
rect 578 -117 585 -115
rect 565 -132 570 -117
rect 580 -132 585 -117
rect 587 -121 595 -104
rect 587 -123 590 -121
rect 592 -123 595 -121
rect 587 -128 595 -123
rect 587 -130 590 -128
rect 592 -130 595 -128
rect 587 -132 595 -130
rect 597 -113 605 -104
rect 597 -115 600 -113
rect 602 -115 605 -113
rect 597 -120 605 -115
rect 597 -122 600 -120
rect 602 -122 605 -120
rect 597 -132 605 -122
rect 607 -121 623 -104
rect 607 -123 612 -121
rect 614 -123 623 -121
rect 607 -128 623 -123
rect 607 -130 612 -128
rect 614 -129 623 -128
rect 625 -129 630 -104
rect 632 -107 637 -104
rect 632 -109 640 -107
rect 632 -111 635 -109
rect 637 -111 640 -109
rect 632 -120 640 -111
rect 642 -120 653 -107
rect 632 -129 637 -120
rect 644 -128 653 -120
rect 614 -130 621 -129
rect 607 -132 621 -130
rect 644 -130 647 -128
rect 649 -130 653 -128
rect 644 -132 653 -130
rect 655 -109 662 -107
rect 655 -111 658 -109
rect 660 -111 662 -109
rect 686 -111 694 -104
rect 655 -116 662 -111
rect 655 -118 658 -116
rect 660 -118 662 -116
rect 655 -120 662 -118
rect 669 -119 674 -111
rect 655 -132 660 -120
rect 667 -121 674 -119
rect 667 -123 669 -121
rect 671 -123 674 -121
rect 667 -125 674 -123
rect 669 -132 674 -125
rect 676 -132 681 -111
rect 683 -122 694 -111
rect 696 -109 701 -104
rect 710 -106 717 -104
rect 710 -108 712 -106
rect 714 -108 717 -106
rect 696 -111 703 -109
rect 710 -110 717 -108
rect 696 -113 699 -111
rect 701 -113 703 -111
rect 712 -112 717 -110
rect 719 -112 725 -104
rect 696 -118 703 -113
rect 696 -120 699 -118
rect 701 -120 703 -118
rect 696 -122 703 -120
rect 721 -116 725 -112
rect 774 -106 781 -104
rect 774 -108 776 -106
rect 778 -108 781 -106
rect 774 -110 781 -108
rect 776 -112 781 -110
rect 783 -112 789 -104
rect 756 -116 761 -114
rect 721 -120 727 -116
rect 683 -128 692 -122
rect 683 -130 688 -128
rect 690 -130 692 -128
rect 720 -128 727 -120
rect 683 -132 692 -130
rect 720 -130 722 -128
rect 724 -130 727 -128
rect 720 -132 727 -130
rect 729 -132 734 -116
rect 736 -118 744 -116
rect 736 -120 739 -118
rect 741 -120 744 -118
rect 736 -132 744 -120
rect 746 -132 751 -116
rect 753 -128 761 -116
rect 753 -130 756 -128
rect 758 -130 761 -128
rect 753 -132 761 -130
rect 763 -119 768 -114
rect 785 -116 789 -112
rect 820 -116 825 -114
rect 763 -121 770 -119
rect 785 -120 791 -116
rect 763 -123 766 -121
rect 768 -123 770 -121
rect 763 -125 770 -123
rect 763 -132 768 -125
rect 784 -128 791 -120
rect 784 -130 786 -128
rect 788 -130 791 -128
rect 784 -132 791 -130
rect 793 -132 798 -116
rect 800 -118 808 -116
rect 800 -120 803 -118
rect 805 -120 808 -118
rect 800 -132 808 -120
rect 810 -132 815 -116
rect 817 -128 825 -116
rect 817 -130 820 -128
rect 822 -130 825 -128
rect 817 -132 825 -130
rect 827 -119 832 -114
rect 827 -121 834 -119
rect 827 -123 830 -121
rect 832 -123 834 -121
rect 827 -125 834 -123
rect 827 -132 832 -125
rect 434 -165 439 -144
rect 432 -167 439 -165
rect 432 -169 434 -167
rect 436 -169 439 -167
rect 432 -171 439 -169
rect 441 -146 453 -144
rect 441 -148 444 -146
rect 446 -148 453 -146
rect 441 -153 453 -148
rect 470 -153 475 -144
rect 441 -155 444 -153
rect 446 -155 455 -153
rect 441 -171 455 -155
rect 457 -160 465 -153
rect 457 -162 460 -160
rect 462 -162 465 -160
rect 457 -167 465 -162
rect 457 -169 460 -167
rect 462 -169 465 -167
rect 457 -171 465 -169
rect 467 -160 475 -153
rect 467 -162 470 -160
rect 472 -162 475 -160
rect 467 -171 475 -162
rect 477 -150 482 -144
rect 477 -152 484 -150
rect 477 -154 480 -152
rect 482 -154 484 -152
rect 477 -156 484 -154
rect 490 -156 495 -144
rect 477 -171 482 -156
rect 488 -158 495 -156
rect 488 -160 490 -158
rect 492 -160 495 -158
rect 488 -165 495 -160
rect 488 -167 490 -165
rect 492 -167 495 -165
rect 488 -169 495 -167
rect 497 -146 506 -144
rect 497 -148 501 -146
rect 503 -148 506 -146
rect 529 -146 543 -144
rect 529 -147 536 -146
rect 497 -156 506 -148
rect 513 -156 518 -147
rect 497 -169 508 -156
rect 510 -165 518 -156
rect 510 -167 513 -165
rect 515 -167 518 -165
rect 510 -169 518 -167
rect 513 -172 518 -169
rect 520 -172 525 -147
rect 527 -148 536 -147
rect 538 -148 543 -146
rect 527 -153 543 -148
rect 527 -155 536 -153
rect 538 -155 543 -153
rect 527 -172 543 -155
rect 545 -154 553 -144
rect 545 -156 548 -154
rect 550 -156 553 -154
rect 545 -161 553 -156
rect 545 -163 548 -161
rect 550 -163 553 -161
rect 545 -172 553 -163
rect 555 -146 563 -144
rect 555 -148 558 -146
rect 560 -148 563 -146
rect 555 -153 563 -148
rect 555 -155 558 -153
rect 560 -155 563 -153
rect 555 -172 563 -155
rect 565 -159 570 -144
rect 580 -159 585 -144
rect 565 -161 572 -159
rect 565 -163 568 -161
rect 570 -163 572 -161
rect 565 -168 572 -163
rect 565 -170 568 -168
rect 570 -170 572 -168
rect 565 -172 572 -170
rect 578 -161 585 -159
rect 578 -163 580 -161
rect 582 -163 585 -161
rect 578 -168 585 -163
rect 578 -170 580 -168
rect 582 -170 585 -168
rect 578 -172 585 -170
rect 587 -146 595 -144
rect 587 -148 590 -146
rect 592 -148 595 -146
rect 587 -153 595 -148
rect 587 -155 590 -153
rect 592 -155 595 -153
rect 587 -172 595 -155
rect 597 -154 605 -144
rect 597 -156 600 -154
rect 602 -156 605 -154
rect 597 -161 605 -156
rect 597 -163 600 -161
rect 602 -163 605 -161
rect 597 -172 605 -163
rect 607 -146 621 -144
rect 607 -148 612 -146
rect 614 -147 621 -146
rect 644 -146 653 -144
rect 614 -148 623 -147
rect 607 -153 623 -148
rect 607 -155 612 -153
rect 614 -155 623 -153
rect 607 -172 623 -155
rect 625 -172 630 -147
rect 632 -156 637 -147
rect 644 -148 647 -146
rect 649 -148 653 -146
rect 644 -156 653 -148
rect 632 -165 640 -156
rect 632 -167 635 -165
rect 637 -167 640 -165
rect 632 -169 640 -167
rect 642 -169 653 -156
rect 655 -156 660 -144
rect 669 -151 674 -144
rect 667 -153 674 -151
rect 667 -155 669 -153
rect 671 -155 674 -153
rect 655 -158 662 -156
rect 667 -157 674 -155
rect 655 -160 658 -158
rect 660 -160 662 -158
rect 655 -165 662 -160
rect 669 -165 674 -157
rect 676 -165 681 -144
rect 683 -146 692 -144
rect 683 -148 688 -146
rect 690 -148 692 -146
rect 720 -146 727 -144
rect 683 -154 692 -148
rect 720 -148 722 -146
rect 724 -148 727 -146
rect 683 -165 694 -154
rect 655 -167 658 -165
rect 660 -167 662 -165
rect 655 -169 662 -167
rect 632 -172 637 -169
rect 686 -172 694 -165
rect 696 -156 703 -154
rect 696 -158 699 -156
rect 701 -158 703 -156
rect 696 -163 703 -158
rect 720 -156 727 -148
rect 696 -165 699 -163
rect 701 -165 703 -163
rect 721 -160 727 -156
rect 729 -160 734 -144
rect 736 -156 744 -144
rect 736 -158 739 -156
rect 741 -158 744 -156
rect 736 -160 744 -158
rect 746 -160 751 -144
rect 753 -146 761 -144
rect 753 -148 756 -146
rect 758 -148 761 -146
rect 753 -160 761 -148
rect 721 -164 725 -160
rect 696 -167 703 -165
rect 712 -166 717 -164
rect 696 -172 701 -167
rect 710 -168 717 -166
rect 710 -170 712 -168
rect 714 -170 717 -168
rect 710 -172 717 -170
rect 719 -172 725 -164
rect 756 -162 761 -160
rect 763 -151 768 -144
rect 784 -146 791 -144
rect 784 -148 786 -146
rect 788 -148 791 -146
rect 763 -153 770 -151
rect 763 -155 766 -153
rect 768 -155 770 -153
rect 763 -157 770 -155
rect 784 -156 791 -148
rect 763 -162 768 -157
rect 785 -160 791 -156
rect 793 -160 798 -144
rect 800 -156 808 -144
rect 800 -158 803 -156
rect 805 -158 808 -156
rect 800 -160 808 -158
rect 810 -160 815 -144
rect 817 -146 825 -144
rect 817 -148 820 -146
rect 822 -148 825 -146
rect 817 -160 825 -148
rect 785 -164 789 -160
rect 776 -166 781 -164
rect 774 -168 781 -166
rect 774 -170 776 -168
rect 778 -170 781 -168
rect 774 -172 781 -170
rect 783 -172 789 -164
rect 820 -162 825 -160
rect 827 -151 832 -144
rect 827 -153 834 -151
rect 827 -155 830 -153
rect 832 -155 834 -153
rect 827 -157 834 -155
rect 827 -162 832 -157
rect 432 -251 439 -249
rect 432 -253 434 -251
rect 436 -253 439 -251
rect 432 -255 439 -253
rect 434 -276 439 -255
rect 441 -265 455 -249
rect 441 -267 444 -265
rect 446 -267 455 -265
rect 457 -251 465 -249
rect 457 -253 460 -251
rect 462 -253 465 -251
rect 457 -258 465 -253
rect 457 -260 460 -258
rect 462 -260 465 -258
rect 457 -267 465 -260
rect 467 -258 475 -249
rect 467 -260 470 -258
rect 472 -260 475 -258
rect 467 -267 475 -260
rect 441 -272 453 -267
rect 441 -274 444 -272
rect 446 -274 453 -272
rect 441 -276 453 -274
rect 470 -276 475 -267
rect 477 -264 482 -249
rect 513 -251 518 -248
rect 488 -253 495 -251
rect 488 -255 490 -253
rect 492 -255 495 -253
rect 488 -260 495 -255
rect 488 -262 490 -260
rect 492 -262 495 -260
rect 488 -264 495 -262
rect 477 -266 484 -264
rect 477 -268 480 -266
rect 482 -268 484 -266
rect 477 -270 484 -268
rect 477 -276 482 -270
rect 490 -276 495 -264
rect 497 -264 508 -251
rect 510 -253 518 -251
rect 510 -255 513 -253
rect 515 -255 518 -253
rect 510 -264 518 -255
rect 497 -272 506 -264
rect 497 -274 501 -272
rect 503 -274 506 -272
rect 513 -273 518 -264
rect 520 -273 525 -248
rect 527 -265 543 -248
rect 527 -267 536 -265
rect 538 -267 543 -265
rect 527 -272 543 -267
rect 527 -273 536 -272
rect 497 -276 506 -274
rect 529 -274 536 -273
rect 538 -274 543 -272
rect 529 -276 543 -274
rect 545 -257 553 -248
rect 545 -259 548 -257
rect 550 -259 553 -257
rect 545 -264 553 -259
rect 545 -266 548 -264
rect 550 -266 553 -264
rect 545 -276 553 -266
rect 555 -265 563 -248
rect 555 -267 558 -265
rect 560 -267 563 -265
rect 555 -272 563 -267
rect 555 -274 558 -272
rect 560 -274 563 -272
rect 555 -276 563 -274
rect 565 -250 572 -248
rect 565 -252 568 -250
rect 570 -252 572 -250
rect 565 -257 572 -252
rect 565 -259 568 -257
rect 570 -259 572 -257
rect 565 -261 572 -259
rect 578 -250 585 -248
rect 578 -252 580 -250
rect 582 -252 585 -250
rect 578 -257 585 -252
rect 578 -259 580 -257
rect 582 -259 585 -257
rect 578 -261 585 -259
rect 565 -276 570 -261
rect 580 -276 585 -261
rect 587 -265 595 -248
rect 587 -267 590 -265
rect 592 -267 595 -265
rect 587 -272 595 -267
rect 587 -274 590 -272
rect 592 -274 595 -272
rect 587 -276 595 -274
rect 597 -257 605 -248
rect 597 -259 600 -257
rect 602 -259 605 -257
rect 597 -264 605 -259
rect 597 -266 600 -264
rect 602 -266 605 -264
rect 597 -276 605 -266
rect 607 -265 623 -248
rect 607 -267 612 -265
rect 614 -267 623 -265
rect 607 -272 623 -267
rect 607 -274 612 -272
rect 614 -273 623 -272
rect 625 -273 630 -248
rect 632 -251 637 -248
rect 632 -253 640 -251
rect 632 -255 635 -253
rect 637 -255 640 -253
rect 632 -264 640 -255
rect 642 -264 653 -251
rect 632 -273 637 -264
rect 644 -272 653 -264
rect 614 -274 621 -273
rect 607 -276 621 -274
rect 644 -274 647 -272
rect 649 -274 653 -272
rect 644 -276 653 -274
rect 655 -253 662 -251
rect 655 -255 658 -253
rect 660 -255 662 -253
rect 686 -255 694 -248
rect 655 -260 662 -255
rect 655 -262 658 -260
rect 660 -262 662 -260
rect 655 -264 662 -262
rect 669 -263 674 -255
rect 655 -276 660 -264
rect 667 -265 674 -263
rect 667 -267 669 -265
rect 671 -267 674 -265
rect 667 -269 674 -267
rect 669 -276 674 -269
rect 676 -276 681 -255
rect 683 -266 694 -255
rect 696 -253 701 -248
rect 710 -250 717 -248
rect 710 -252 712 -250
rect 714 -252 717 -250
rect 696 -255 703 -253
rect 710 -254 717 -252
rect 696 -257 699 -255
rect 701 -257 703 -255
rect 712 -256 717 -254
rect 719 -256 725 -248
rect 696 -262 703 -257
rect 696 -264 699 -262
rect 701 -264 703 -262
rect 696 -266 703 -264
rect 721 -260 725 -256
rect 774 -250 781 -248
rect 774 -252 776 -250
rect 778 -252 781 -250
rect 774 -254 781 -252
rect 776 -256 781 -254
rect 783 -256 789 -248
rect 756 -260 761 -258
rect 721 -264 727 -260
rect 683 -272 692 -266
rect 683 -274 688 -272
rect 690 -274 692 -272
rect 720 -272 727 -264
rect 683 -276 692 -274
rect 720 -274 722 -272
rect 724 -274 727 -272
rect 720 -276 727 -274
rect 729 -276 734 -260
rect 736 -262 744 -260
rect 736 -264 739 -262
rect 741 -264 744 -262
rect 736 -276 744 -264
rect 746 -276 751 -260
rect 753 -272 761 -260
rect 753 -274 756 -272
rect 758 -274 761 -272
rect 753 -276 761 -274
rect 763 -263 768 -258
rect 785 -260 789 -256
rect 820 -260 825 -258
rect 763 -265 770 -263
rect 785 -264 791 -260
rect 763 -267 766 -265
rect 768 -267 770 -265
rect 763 -269 770 -267
rect 763 -276 768 -269
rect 784 -272 791 -264
rect 784 -274 786 -272
rect 788 -274 791 -272
rect 784 -276 791 -274
rect 793 -276 798 -260
rect 800 -262 808 -260
rect 800 -264 803 -262
rect 805 -264 808 -262
rect 800 -276 808 -264
rect 810 -276 815 -260
rect 817 -272 825 -260
rect 817 -274 820 -272
rect 822 -274 825 -272
rect 817 -276 825 -274
rect 827 -263 832 -258
rect 827 -265 834 -263
rect 827 -267 830 -265
rect 832 -267 834 -265
rect 827 -269 834 -267
rect 827 -276 832 -269
<< alu1 >>
rect 2 293 838 294
rect 2 291 26 293
rect 28 291 159 293
rect 161 291 399 293
rect 401 291 584 293
rect 586 291 776 293
rect 778 291 838 293
rect 2 289 838 291
rect 2 287 37 289
rect 39 287 77 289
rect 79 287 296 289
rect 298 287 344 289
rect 346 287 563 289
rect 565 287 611 289
rect 613 287 830 289
rect 832 287 838 289
rect 2 286 838 287
rect 6 266 10 273
rect 37 272 42 274
rect 6 264 7 266
rect 9 264 10 266
rect 6 263 19 264
rect 6 261 11 263
rect 13 261 19 263
rect 6 260 19 261
rect 13 255 27 256
rect 13 253 21 255
rect 23 253 27 255
rect 13 252 27 253
rect 37 270 38 272
rect 40 270 42 272
rect 37 265 42 270
rect 37 263 38 265
rect 40 263 42 265
rect 37 261 42 263
rect 13 246 18 252
rect 13 244 15 246
rect 17 244 18 246
rect 13 243 18 244
rect 38 260 42 261
rect 46 272 50 273
rect 46 270 47 272
rect 49 270 50 272
rect 46 264 50 270
rect 297 280 301 281
rect 288 276 301 280
rect 86 274 91 276
rect 77 272 82 274
rect 46 263 59 264
rect 46 261 51 263
rect 53 261 59 263
rect 46 260 59 261
rect 38 258 39 260
rect 41 258 42 260
rect 38 241 42 258
rect 53 255 67 256
rect 53 253 61 255
rect 63 253 67 255
rect 53 252 67 253
rect 77 270 78 272
rect 80 270 82 272
rect 77 265 82 270
rect 77 263 78 265
rect 80 263 82 265
rect 77 261 82 263
rect 53 249 58 252
rect 53 247 55 249
rect 57 247 58 249
rect 53 243 58 247
rect 78 255 82 261
rect 78 253 79 255
rect 81 253 82 255
rect 30 239 38 241
rect 40 239 42 241
rect 78 241 82 253
rect 30 235 42 239
rect 70 239 78 241
rect 80 239 82 241
rect 70 235 82 239
rect 86 272 88 274
rect 90 272 91 274
rect 86 267 91 272
rect 86 265 88 267
rect 90 265 91 267
rect 86 263 91 265
rect 86 247 90 263
rect 117 263 155 264
rect 117 261 119 263
rect 121 261 155 263
rect 117 260 155 261
rect 117 257 122 260
rect 114 255 122 257
rect 114 253 115 255
rect 117 253 122 255
rect 114 251 122 253
rect 132 255 147 256
rect 132 253 134 255
rect 136 253 137 255
rect 139 253 141 255
rect 143 253 147 255
rect 132 252 147 253
rect 86 245 87 247
rect 89 245 90 247
rect 86 241 90 245
rect 86 239 91 241
rect 134 243 138 252
rect 165 271 171 273
rect 165 269 166 271
rect 168 269 171 271
rect 165 264 171 269
rect 165 262 166 264
rect 168 262 171 264
rect 165 260 171 262
rect 167 255 171 260
rect 167 253 168 255
rect 170 253 171 255
rect 167 240 171 253
rect 86 237 88 239
rect 90 237 91 239
rect 86 235 91 237
rect 165 239 171 240
rect 165 237 166 239
rect 168 237 171 239
rect 165 236 171 237
rect 175 271 181 273
rect 255 274 260 276
rect 255 272 256 274
rect 258 272 260 274
rect 175 269 178 271
rect 180 269 181 271
rect 175 268 181 269
rect 175 266 178 268
rect 180 266 181 268
rect 175 264 181 266
rect 175 262 178 264
rect 180 262 181 264
rect 175 260 181 262
rect 175 240 179 260
rect 191 263 229 264
rect 191 261 208 263
rect 210 261 229 263
rect 191 260 229 261
rect 224 257 229 260
rect 199 255 214 256
rect 199 253 203 255
rect 205 253 210 255
rect 212 253 214 255
rect 199 252 214 253
rect 224 255 232 257
rect 224 253 229 255
rect 231 253 232 255
rect 208 247 212 252
rect 224 251 232 253
rect 255 267 260 272
rect 255 265 256 267
rect 258 265 260 267
rect 255 263 260 265
rect 208 245 209 247
rect 211 245 212 247
rect 208 243 212 245
rect 175 239 181 240
rect 175 237 178 239
rect 180 237 181 239
rect 175 236 181 237
rect 256 244 260 263
rect 265 272 269 273
rect 265 270 266 272
rect 268 270 269 272
rect 265 264 269 270
rect 265 262 286 264
rect 265 260 270 262
rect 272 260 286 262
rect 256 242 257 244
rect 259 242 260 244
rect 265 255 286 256
rect 265 253 266 255
rect 268 253 280 255
rect 282 253 286 255
rect 265 252 286 253
rect 299 274 301 276
rect 297 269 301 274
rect 299 267 301 269
rect 265 243 269 252
rect 297 251 301 267
rect 313 272 317 273
rect 313 270 314 272
rect 316 270 317 272
rect 313 264 317 270
rect 564 280 568 281
rect 555 276 568 280
rect 353 274 358 276
rect 344 272 349 274
rect 313 263 326 264
rect 313 261 318 263
rect 320 261 326 263
rect 313 260 326 261
rect 297 249 298 251
rect 300 249 301 251
rect 297 248 301 249
rect 296 246 301 248
rect 296 244 297 246
rect 299 244 301 246
rect 296 242 301 244
rect 320 255 334 256
rect 320 253 328 255
rect 330 253 334 255
rect 320 252 334 253
rect 344 270 345 272
rect 347 270 349 272
rect 344 265 349 270
rect 344 263 345 265
rect 347 263 349 265
rect 344 261 349 263
rect 320 249 325 252
rect 320 247 322 249
rect 324 247 325 249
rect 320 243 325 247
rect 345 255 349 261
rect 345 253 346 255
rect 348 253 349 255
rect 256 241 260 242
rect 255 239 260 241
rect 345 241 349 253
rect 255 237 256 239
rect 258 237 260 239
rect 255 235 260 237
rect 337 239 345 241
rect 347 239 349 241
rect 337 235 349 239
rect 353 272 355 274
rect 357 272 358 274
rect 353 267 358 272
rect 353 265 355 267
rect 357 265 358 267
rect 353 263 358 265
rect 353 247 357 263
rect 384 263 422 264
rect 384 261 386 263
rect 388 261 422 263
rect 384 260 422 261
rect 384 257 389 260
rect 381 255 389 257
rect 381 253 382 255
rect 384 253 389 255
rect 381 251 389 253
rect 399 255 414 256
rect 399 253 401 255
rect 403 253 404 255
rect 406 253 408 255
rect 410 253 414 255
rect 399 252 414 253
rect 353 245 354 247
rect 356 245 357 247
rect 353 241 357 245
rect 353 239 358 241
rect 401 243 405 252
rect 432 271 438 273
rect 432 269 433 271
rect 435 269 438 271
rect 432 264 438 269
rect 432 262 433 264
rect 435 262 438 264
rect 432 260 438 262
rect 434 255 438 260
rect 434 253 435 255
rect 437 253 438 255
rect 434 240 438 253
rect 353 237 355 239
rect 357 237 358 239
rect 353 235 358 237
rect 432 239 438 240
rect 432 237 433 239
rect 435 237 438 239
rect 432 236 438 237
rect 442 271 448 273
rect 522 274 527 276
rect 522 272 523 274
rect 525 272 527 274
rect 442 269 445 271
rect 447 269 448 271
rect 442 268 448 269
rect 442 266 445 268
rect 447 266 448 268
rect 442 264 448 266
rect 442 262 445 264
rect 447 262 448 264
rect 442 260 448 262
rect 442 240 446 260
rect 458 263 496 264
rect 458 261 475 263
rect 477 261 496 263
rect 458 260 496 261
rect 491 257 496 260
rect 466 255 481 256
rect 466 253 470 255
rect 472 253 477 255
rect 479 253 481 255
rect 466 252 481 253
rect 491 255 499 257
rect 491 253 496 255
rect 498 253 499 255
rect 475 247 479 252
rect 491 251 499 253
rect 522 267 527 272
rect 522 265 523 267
rect 525 265 527 267
rect 522 263 527 265
rect 475 245 476 247
rect 478 245 479 247
rect 475 243 479 245
rect 442 239 448 240
rect 442 237 445 239
rect 447 237 448 239
rect 442 236 448 237
rect 523 245 527 263
rect 532 272 536 273
rect 532 270 533 272
rect 535 270 536 272
rect 532 264 536 270
rect 532 262 553 264
rect 532 260 537 262
rect 539 260 553 262
rect 523 243 524 245
rect 526 243 527 245
rect 532 255 553 256
rect 532 253 533 255
rect 535 253 547 255
rect 549 253 553 255
rect 532 252 553 253
rect 566 274 568 276
rect 564 269 568 274
rect 566 267 568 269
rect 532 243 536 252
rect 564 251 568 267
rect 580 272 584 273
rect 580 270 581 272
rect 583 270 584 272
rect 580 264 584 270
rect 831 280 835 281
rect 822 276 835 280
rect 620 274 625 276
rect 611 272 616 274
rect 580 263 593 264
rect 580 261 585 263
rect 587 261 593 263
rect 580 260 593 261
rect 564 249 565 251
rect 567 249 568 251
rect 564 248 568 249
rect 563 246 568 248
rect 563 244 564 246
rect 566 244 568 246
rect 523 241 527 243
rect 563 242 568 244
rect 587 255 601 256
rect 587 253 595 255
rect 597 253 601 255
rect 587 252 601 253
rect 611 270 612 272
rect 614 270 616 272
rect 611 265 616 270
rect 611 263 612 265
rect 614 263 616 265
rect 611 261 616 263
rect 587 249 592 252
rect 587 247 589 249
rect 591 247 592 249
rect 587 243 592 247
rect 612 255 616 261
rect 612 253 613 255
rect 615 253 616 255
rect 522 239 527 241
rect 612 241 616 253
rect 522 237 523 239
rect 525 237 527 239
rect 522 235 527 237
rect 604 239 612 241
rect 614 239 616 241
rect 604 235 616 239
rect 620 272 622 274
rect 624 272 625 274
rect 620 267 625 272
rect 620 265 622 267
rect 624 265 625 267
rect 620 263 625 265
rect 620 247 624 263
rect 651 263 689 264
rect 651 261 653 263
rect 655 261 689 263
rect 651 260 689 261
rect 651 257 656 260
rect 648 255 656 257
rect 648 253 649 255
rect 651 253 656 255
rect 648 251 656 253
rect 666 255 681 256
rect 666 253 668 255
rect 670 253 671 255
rect 673 253 675 255
rect 677 253 681 255
rect 666 252 681 253
rect 620 245 621 247
rect 623 245 624 247
rect 620 241 624 245
rect 620 239 625 241
rect 668 243 672 252
rect 699 271 705 273
rect 699 269 700 271
rect 702 269 705 271
rect 699 264 705 269
rect 699 262 700 264
rect 702 262 705 264
rect 699 260 705 262
rect 701 255 705 260
rect 701 253 702 255
rect 704 253 705 255
rect 701 240 705 253
rect 620 237 622 239
rect 624 237 625 239
rect 620 235 625 237
rect 699 239 705 240
rect 699 237 700 239
rect 702 237 705 239
rect 699 236 705 237
rect 709 271 715 273
rect 789 274 794 276
rect 789 272 790 274
rect 792 272 794 274
rect 709 269 712 271
rect 714 269 715 271
rect 709 268 715 269
rect 709 266 712 268
rect 714 266 715 268
rect 709 264 715 266
rect 709 262 712 264
rect 714 262 715 264
rect 709 260 715 262
rect 709 240 713 260
rect 725 263 763 264
rect 725 261 742 263
rect 744 261 763 263
rect 725 260 763 261
rect 758 257 763 260
rect 733 255 748 256
rect 733 253 737 255
rect 739 253 744 255
rect 746 253 748 255
rect 733 252 748 253
rect 758 255 766 257
rect 758 253 763 255
rect 765 253 766 255
rect 742 247 746 252
rect 758 251 766 253
rect 789 267 794 272
rect 789 265 790 267
rect 792 265 794 267
rect 789 263 794 265
rect 742 245 743 247
rect 745 245 746 247
rect 742 243 746 245
rect 709 239 715 240
rect 709 237 712 239
rect 714 237 715 239
rect 709 236 715 237
rect 790 245 794 263
rect 799 272 803 273
rect 799 270 800 272
rect 802 270 803 272
rect 799 264 803 270
rect 799 262 820 264
rect 799 260 804 262
rect 806 260 820 262
rect 790 243 791 245
rect 793 243 794 245
rect 799 255 820 256
rect 799 253 800 255
rect 802 253 814 255
rect 816 253 820 255
rect 799 252 820 253
rect 833 274 835 276
rect 831 269 835 274
rect 833 267 835 269
rect 799 243 803 252
rect 831 251 835 267
rect 831 249 832 251
rect 834 249 835 251
rect 831 248 835 249
rect 830 246 835 248
rect 830 244 831 246
rect 833 244 835 246
rect 790 241 794 243
rect 830 242 835 244
rect 789 239 794 241
rect 789 237 790 239
rect 792 237 794 239
rect 789 235 794 237
rect 2 229 838 230
rect 2 227 27 229
rect 29 227 37 229
rect 39 227 67 229
rect 69 227 77 229
rect 79 227 296 229
rect 298 227 334 229
rect 336 227 344 229
rect 346 227 563 229
rect 565 227 601 229
rect 603 227 611 229
rect 613 227 830 229
rect 832 227 838 229
rect 2 226 838 227
rect 2 224 214 226
rect 216 224 481 226
rect 483 224 748 226
rect 750 224 838 226
rect 2 223 838 224
rect 2 221 769 223
rect 771 221 838 223
rect 2 217 838 221
rect 2 215 27 217
rect 29 215 37 217
rect 39 215 67 217
rect 69 215 77 217
rect 79 215 296 217
rect 298 215 334 217
rect 336 215 344 217
rect 346 215 563 217
rect 565 215 601 217
rect 603 215 611 217
rect 613 215 830 217
rect 832 215 838 217
rect 2 214 838 215
rect 13 195 18 201
rect 30 205 42 209
rect 30 203 38 205
rect 40 203 42 205
rect 13 193 15 195
rect 17 193 18 195
rect 13 192 18 193
rect 13 191 27 192
rect 13 189 21 191
rect 23 189 27 191
rect 13 188 27 189
rect 6 183 19 184
rect 6 181 11 183
rect 13 181 19 183
rect 6 180 19 181
rect 6 174 10 180
rect 38 183 42 203
rect 53 197 58 201
rect 53 195 55 197
rect 57 195 58 197
rect 70 205 82 209
rect 70 203 78 205
rect 80 203 82 205
rect 53 192 58 195
rect 53 191 67 192
rect 53 189 61 191
rect 63 189 67 191
rect 53 188 67 189
rect 6 172 7 174
rect 9 172 10 174
rect 6 171 10 172
rect 37 181 39 183
rect 41 181 42 183
rect 37 180 42 181
rect 37 178 38 180
rect 40 178 42 180
rect 37 172 42 178
rect 37 170 38 172
rect 40 170 42 172
rect 46 183 59 184
rect 46 181 51 183
rect 53 181 59 183
rect 46 180 59 181
rect 46 175 50 180
rect 78 191 82 203
rect 78 189 79 191
rect 81 189 82 191
rect 78 183 82 189
rect 46 173 47 175
rect 49 173 50 175
rect 46 171 50 173
rect 77 181 82 183
rect 77 179 78 181
rect 80 179 82 181
rect 77 174 82 179
rect 37 168 42 170
rect 77 172 78 174
rect 80 172 82 174
rect 77 170 82 172
rect 86 207 91 209
rect 86 205 88 207
rect 90 205 91 207
rect 86 203 91 205
rect 86 199 90 203
rect 86 197 87 199
rect 89 197 90 199
rect 86 181 90 197
rect 165 207 171 208
rect 165 205 166 207
rect 168 205 171 207
rect 165 204 171 205
rect 86 179 91 181
rect 86 177 88 179
rect 90 177 91 179
rect 86 172 91 177
rect 114 191 122 193
rect 134 192 138 201
rect 114 189 115 191
rect 117 189 122 191
rect 114 187 122 189
rect 132 191 147 192
rect 132 189 134 191
rect 136 189 137 191
rect 139 189 141 191
rect 143 189 147 191
rect 132 188 147 189
rect 117 184 122 187
rect 167 191 171 204
rect 167 189 168 191
rect 170 189 171 191
rect 117 183 155 184
rect 117 181 132 183
rect 134 181 155 183
rect 117 180 155 181
rect 167 184 171 189
rect 165 182 171 184
rect 165 180 166 182
rect 168 180 171 182
rect 165 175 171 180
rect 165 173 166 175
rect 168 173 171 175
rect 86 170 88 172
rect 90 170 91 172
rect 86 168 91 170
rect 165 171 171 173
rect 175 207 181 208
rect 175 205 178 207
rect 180 205 181 207
rect 175 204 181 205
rect 255 207 262 209
rect 255 205 256 207
rect 258 205 259 207
rect 261 205 262 207
rect 175 184 179 204
rect 208 199 212 201
rect 208 197 209 199
rect 211 197 212 199
rect 175 182 181 184
rect 175 180 178 182
rect 180 180 181 182
rect 175 178 181 180
rect 175 176 178 178
rect 180 176 181 178
rect 175 175 181 176
rect 175 173 178 175
rect 180 173 181 175
rect 175 171 181 173
rect 208 192 212 197
rect 255 203 262 205
rect 199 191 214 192
rect 199 189 203 191
rect 205 189 210 191
rect 212 189 214 191
rect 199 188 214 189
rect 224 191 232 193
rect 224 189 229 191
rect 231 189 232 191
rect 224 187 232 189
rect 224 186 229 187
rect 224 184 226 186
rect 228 184 229 186
rect 191 180 229 184
rect 256 181 260 203
rect 265 197 269 198
rect 265 195 266 197
rect 268 195 269 197
rect 265 192 269 195
rect 265 191 286 192
rect 265 189 280 191
rect 282 189 286 191
rect 265 188 286 189
rect 296 200 301 202
rect 296 198 297 200
rect 299 198 301 200
rect 296 196 301 198
rect 255 179 260 181
rect 255 177 256 179
rect 258 177 260 179
rect 255 172 260 177
rect 255 170 256 172
rect 258 170 260 172
rect 265 182 270 184
rect 272 182 286 184
rect 265 180 286 182
rect 265 178 269 180
rect 265 176 266 178
rect 268 176 269 178
rect 265 171 269 176
rect 255 168 260 170
rect 297 177 301 196
rect 320 198 325 201
rect 320 196 322 198
rect 324 196 325 198
rect 337 205 349 209
rect 337 203 345 205
rect 347 203 349 205
rect 320 192 325 196
rect 320 191 334 192
rect 320 189 328 191
rect 330 189 334 191
rect 320 188 334 189
rect 299 175 301 177
rect 297 170 301 175
rect 313 183 326 184
rect 313 181 318 183
rect 320 181 326 183
rect 313 180 326 181
rect 313 175 317 180
rect 345 191 349 203
rect 345 189 346 191
rect 348 189 349 191
rect 345 183 349 189
rect 313 173 314 175
rect 316 173 317 175
rect 313 171 317 173
rect 344 181 349 183
rect 344 179 345 181
rect 347 179 349 181
rect 344 174 349 179
rect 299 168 301 170
rect 288 167 301 168
rect 288 165 290 167
rect 292 165 301 167
rect 288 164 301 165
rect 297 163 301 164
rect 344 172 345 174
rect 347 172 349 174
rect 344 170 349 172
rect 353 207 358 209
rect 353 205 355 207
rect 357 205 358 207
rect 353 203 358 205
rect 353 199 357 203
rect 353 197 354 199
rect 356 197 357 199
rect 353 181 357 197
rect 432 207 438 208
rect 432 205 433 207
rect 435 205 438 207
rect 432 204 438 205
rect 353 179 358 181
rect 353 177 355 179
rect 357 177 358 179
rect 353 172 358 177
rect 381 191 389 193
rect 401 192 405 201
rect 381 189 382 191
rect 384 189 389 191
rect 381 187 389 189
rect 399 191 414 192
rect 399 189 401 191
rect 403 189 404 191
rect 406 189 408 191
rect 410 189 414 191
rect 399 188 414 189
rect 384 184 389 187
rect 434 191 438 204
rect 434 189 435 191
rect 437 189 438 191
rect 384 183 422 184
rect 384 181 399 183
rect 401 181 422 183
rect 384 180 422 181
rect 434 184 438 189
rect 432 182 438 184
rect 432 180 433 182
rect 435 180 438 182
rect 432 175 438 180
rect 432 173 433 175
rect 435 173 438 175
rect 353 170 355 172
rect 357 170 358 172
rect 353 168 358 170
rect 432 171 438 173
rect 442 207 448 208
rect 442 205 445 207
rect 447 205 448 207
rect 442 204 448 205
rect 522 207 529 209
rect 522 205 523 207
rect 525 205 526 207
rect 528 205 529 207
rect 442 184 446 204
rect 475 199 479 201
rect 475 197 476 199
rect 478 197 479 199
rect 442 182 448 184
rect 442 180 445 182
rect 447 180 448 182
rect 442 178 448 180
rect 442 176 445 178
rect 447 176 448 178
rect 442 175 448 176
rect 442 173 445 175
rect 447 173 448 175
rect 442 171 448 173
rect 475 192 479 197
rect 522 203 529 205
rect 466 191 481 192
rect 466 189 470 191
rect 472 189 477 191
rect 479 189 481 191
rect 466 188 481 189
rect 491 191 499 193
rect 491 189 496 191
rect 498 189 499 191
rect 491 187 499 189
rect 491 186 496 187
rect 491 184 493 186
rect 495 184 496 186
rect 458 180 496 184
rect 523 181 527 203
rect 532 197 536 198
rect 532 195 533 197
rect 535 195 536 197
rect 532 192 536 195
rect 532 191 553 192
rect 532 189 547 191
rect 549 189 553 191
rect 532 188 553 189
rect 563 200 568 202
rect 563 198 564 200
rect 566 198 568 200
rect 563 196 568 198
rect 522 179 527 181
rect 522 177 523 179
rect 525 177 527 179
rect 522 172 527 177
rect 522 170 523 172
rect 525 170 527 172
rect 532 182 537 184
rect 539 182 553 184
rect 532 180 553 182
rect 532 178 536 180
rect 532 176 533 178
rect 535 176 536 178
rect 532 171 536 176
rect 522 168 527 170
rect 564 177 568 196
rect 587 196 592 201
rect 604 205 616 209
rect 604 203 612 205
rect 614 203 616 205
rect 587 194 588 196
rect 590 194 592 196
rect 587 192 592 194
rect 587 191 601 192
rect 587 189 595 191
rect 597 189 601 191
rect 587 188 601 189
rect 566 175 568 177
rect 564 170 568 175
rect 580 183 593 184
rect 580 181 585 183
rect 587 181 593 183
rect 580 180 593 181
rect 580 175 584 180
rect 612 191 616 203
rect 612 189 613 191
rect 615 189 616 191
rect 612 183 616 189
rect 580 173 581 175
rect 583 173 584 175
rect 580 171 584 173
rect 611 181 616 183
rect 611 179 612 181
rect 614 179 616 181
rect 611 174 616 179
rect 566 168 568 170
rect 555 167 568 168
rect 555 165 557 167
rect 559 165 568 167
rect 555 164 568 165
rect 564 163 568 164
rect 611 172 612 174
rect 614 172 616 174
rect 611 170 616 172
rect 620 207 625 209
rect 620 205 622 207
rect 624 205 625 207
rect 620 203 625 205
rect 620 199 624 203
rect 620 197 621 199
rect 623 197 624 199
rect 620 181 624 197
rect 699 207 705 208
rect 699 205 700 207
rect 702 205 705 207
rect 699 204 705 205
rect 620 179 625 181
rect 620 177 622 179
rect 624 177 625 179
rect 620 172 625 177
rect 648 191 656 193
rect 668 192 672 201
rect 648 189 649 191
rect 651 189 656 191
rect 648 187 656 189
rect 666 191 681 192
rect 666 189 668 191
rect 670 189 671 191
rect 673 189 675 191
rect 677 189 681 191
rect 666 188 681 189
rect 651 184 656 187
rect 701 191 705 204
rect 701 189 702 191
rect 704 189 705 191
rect 651 183 689 184
rect 651 181 666 183
rect 668 181 689 183
rect 651 180 689 181
rect 701 184 705 189
rect 699 182 705 184
rect 699 180 700 182
rect 702 180 705 182
rect 699 175 705 180
rect 699 173 700 175
rect 702 173 705 175
rect 620 170 622 172
rect 624 170 625 172
rect 620 168 625 170
rect 699 171 705 173
rect 709 207 715 208
rect 709 205 712 207
rect 714 205 715 207
rect 709 204 715 205
rect 789 208 796 209
rect 789 207 793 208
rect 789 205 790 207
rect 792 206 793 207
rect 795 206 796 208
rect 792 205 796 206
rect 709 184 713 204
rect 742 199 746 201
rect 742 197 743 199
rect 745 197 746 199
rect 709 182 715 184
rect 709 180 712 182
rect 714 180 715 182
rect 709 178 715 180
rect 709 176 712 178
rect 714 176 715 178
rect 709 175 715 176
rect 709 173 712 175
rect 714 173 715 175
rect 709 171 715 173
rect 742 192 746 197
rect 789 203 796 205
rect 733 191 748 192
rect 733 189 737 191
rect 739 189 744 191
rect 746 189 748 191
rect 733 188 748 189
rect 758 191 766 193
rect 758 189 763 191
rect 765 189 766 191
rect 758 187 766 189
rect 758 186 763 187
rect 758 184 760 186
rect 762 184 763 186
rect 725 180 763 184
rect 790 181 794 203
rect 799 197 803 198
rect 799 195 800 197
rect 802 195 803 197
rect 799 192 803 195
rect 799 191 820 192
rect 799 189 814 191
rect 816 189 820 191
rect 799 188 820 189
rect 830 200 835 202
rect 830 198 831 200
rect 833 198 835 200
rect 830 196 835 198
rect 789 179 794 181
rect 789 177 790 179
rect 792 177 794 179
rect 789 172 794 177
rect 789 170 790 172
rect 792 170 794 172
rect 799 182 804 184
rect 806 182 820 184
rect 799 180 820 182
rect 799 178 803 180
rect 799 176 800 178
rect 802 176 803 178
rect 799 171 803 176
rect 789 168 794 170
rect 831 177 835 196
rect 833 175 835 177
rect 831 170 835 175
rect 833 168 835 170
rect 822 167 835 168
rect 822 165 824 167
rect 826 165 835 167
rect 822 164 835 165
rect 831 163 835 164
rect 2 157 838 158
rect 2 155 37 157
rect 39 155 77 157
rect 79 155 296 157
rect 298 155 344 157
rect 346 155 563 157
rect 565 155 611 157
rect 613 155 830 157
rect 832 155 838 157
rect 2 149 838 155
rect 2 147 833 149
rect 835 147 838 149
rect 2 145 838 147
rect 2 143 8 145
rect 10 143 37 145
rect 39 143 77 145
rect 79 143 296 145
rect 298 143 344 145
rect 346 143 563 145
rect 565 143 611 145
rect 613 143 830 145
rect 832 143 838 145
rect 2 142 838 143
rect 6 122 10 129
rect 37 131 42 133
rect 37 129 38 131
rect 40 129 42 131
rect 6 120 7 122
rect 9 120 10 122
rect 6 119 19 120
rect 6 117 11 119
rect 13 117 19 119
rect 6 116 19 117
rect 13 111 27 112
rect 13 109 21 111
rect 23 109 27 111
rect 13 108 27 109
rect 37 123 42 129
rect 37 121 38 123
rect 40 121 42 123
rect 37 119 42 121
rect 37 117 39 119
rect 41 117 42 119
rect 37 115 42 117
rect 46 128 50 129
rect 46 126 47 128
rect 49 126 50 128
rect 46 120 50 126
rect 297 136 301 137
rect 288 132 301 136
rect 86 130 91 132
rect 77 128 82 130
rect 46 119 59 120
rect 46 117 51 119
rect 53 117 59 119
rect 46 116 59 117
rect 13 103 18 108
rect 13 101 14 103
rect 16 101 18 103
rect 13 100 18 101
rect 38 97 42 115
rect 53 111 67 112
rect 53 109 61 111
rect 63 109 67 111
rect 53 108 67 109
rect 77 126 78 128
rect 80 126 82 128
rect 77 121 82 126
rect 77 119 78 121
rect 80 119 82 121
rect 77 117 82 119
rect 53 106 58 108
rect 53 104 55 106
rect 57 104 58 106
rect 53 99 58 104
rect 78 111 82 117
rect 78 109 79 111
rect 81 109 82 111
rect 30 95 38 97
rect 40 95 42 97
rect 78 97 82 109
rect 30 91 42 95
rect 70 95 78 97
rect 80 95 82 97
rect 70 91 82 95
rect 86 128 88 130
rect 90 128 91 130
rect 86 123 91 128
rect 86 121 88 123
rect 90 121 91 123
rect 86 119 91 121
rect 86 103 90 119
rect 117 119 155 120
rect 117 117 136 119
rect 138 117 155 119
rect 117 116 155 117
rect 117 113 122 116
rect 114 111 122 113
rect 114 109 115 111
rect 117 109 122 111
rect 114 107 122 109
rect 132 111 147 112
rect 132 109 134 111
rect 136 109 138 111
rect 140 109 141 111
rect 143 109 147 111
rect 132 108 147 109
rect 86 101 87 103
rect 89 101 90 103
rect 86 97 90 101
rect 86 95 91 97
rect 134 99 138 108
rect 165 127 171 129
rect 165 125 166 127
rect 168 125 171 127
rect 165 120 171 125
rect 165 118 166 120
rect 168 118 171 120
rect 165 116 171 118
rect 167 111 171 116
rect 167 109 168 111
rect 170 109 171 111
rect 167 96 171 109
rect 86 93 88 95
rect 90 93 91 95
rect 86 91 91 93
rect 165 95 171 96
rect 165 93 166 95
rect 168 93 171 95
rect 165 92 171 93
rect 175 127 181 129
rect 255 130 260 132
rect 255 128 256 130
rect 258 128 260 130
rect 175 125 178 127
rect 180 125 181 127
rect 175 124 181 125
rect 175 122 178 124
rect 180 122 181 124
rect 175 120 181 122
rect 175 118 178 120
rect 180 118 181 120
rect 175 116 181 118
rect 175 96 179 116
rect 191 119 229 120
rect 191 117 226 119
rect 228 117 229 119
rect 191 116 229 117
rect 224 113 229 116
rect 199 111 214 112
rect 199 109 203 111
rect 205 109 210 111
rect 212 109 214 111
rect 199 108 214 109
rect 224 111 232 113
rect 224 109 229 111
rect 231 109 232 111
rect 208 103 212 108
rect 224 107 232 109
rect 255 123 260 128
rect 255 121 256 123
rect 258 121 260 123
rect 255 119 260 121
rect 208 101 209 103
rect 211 101 212 103
rect 208 99 212 101
rect 175 95 181 96
rect 175 93 178 95
rect 180 93 181 95
rect 175 92 181 93
rect 256 97 260 119
rect 265 128 269 129
rect 265 126 266 128
rect 268 126 269 128
rect 265 120 269 126
rect 265 118 286 120
rect 265 116 270 118
rect 272 116 286 118
rect 265 111 286 112
rect 265 109 266 111
rect 268 109 280 111
rect 282 109 286 111
rect 265 108 286 109
rect 299 130 301 132
rect 297 125 301 130
rect 299 123 301 125
rect 265 104 269 108
rect 297 107 301 123
rect 313 124 317 129
rect 313 122 314 124
rect 316 122 317 124
rect 564 136 568 137
rect 555 132 568 136
rect 353 130 358 132
rect 344 128 349 130
rect 313 120 317 122
rect 313 119 326 120
rect 313 117 318 119
rect 320 117 326 119
rect 313 116 326 117
rect 297 105 298 107
rect 300 105 301 107
rect 297 104 301 105
rect 296 102 301 104
rect 296 100 297 102
rect 299 100 301 102
rect 296 98 301 100
rect 320 111 334 112
rect 320 109 328 111
rect 330 109 334 111
rect 320 108 334 109
rect 344 126 345 128
rect 347 126 349 128
rect 344 121 349 126
rect 344 119 345 121
rect 347 119 349 121
rect 344 117 349 119
rect 320 106 325 108
rect 320 104 322 106
rect 324 104 325 106
rect 320 99 325 104
rect 345 111 349 117
rect 345 109 346 111
rect 348 109 349 111
rect 255 95 262 97
rect 345 97 349 109
rect 255 93 256 95
rect 258 93 259 95
rect 261 93 262 95
rect 255 91 262 93
rect 337 95 345 97
rect 347 95 349 97
rect 337 91 349 95
rect 353 128 355 130
rect 357 128 358 130
rect 353 123 358 128
rect 353 121 355 123
rect 357 121 358 123
rect 353 119 358 121
rect 353 103 357 119
rect 384 119 422 120
rect 384 117 403 119
rect 405 117 422 119
rect 384 116 422 117
rect 384 113 389 116
rect 381 111 389 113
rect 381 109 382 111
rect 384 109 389 111
rect 381 107 389 109
rect 399 111 414 112
rect 399 109 401 111
rect 403 109 405 111
rect 407 109 408 111
rect 410 109 414 111
rect 399 108 414 109
rect 353 101 354 103
rect 356 101 357 103
rect 353 97 357 101
rect 353 95 358 97
rect 401 99 405 108
rect 432 127 438 129
rect 432 125 433 127
rect 435 125 438 127
rect 432 120 438 125
rect 432 118 433 120
rect 435 118 438 120
rect 432 116 438 118
rect 434 111 438 116
rect 434 109 435 111
rect 437 109 438 111
rect 434 96 438 109
rect 353 93 355 95
rect 357 93 358 95
rect 353 91 358 93
rect 432 95 438 96
rect 432 93 433 95
rect 435 93 438 95
rect 432 92 438 93
rect 442 127 448 129
rect 522 130 527 132
rect 522 128 523 130
rect 525 128 527 130
rect 442 125 445 127
rect 447 125 448 127
rect 442 124 448 125
rect 442 122 445 124
rect 447 122 448 124
rect 442 120 448 122
rect 442 118 445 120
rect 447 118 448 120
rect 442 116 448 118
rect 442 96 446 116
rect 458 119 496 120
rect 458 117 493 119
rect 495 117 496 119
rect 458 116 496 117
rect 491 113 496 116
rect 466 111 481 112
rect 466 109 470 111
rect 472 109 477 111
rect 479 109 481 111
rect 466 108 481 109
rect 491 111 499 113
rect 491 109 496 111
rect 498 109 499 111
rect 475 103 479 108
rect 491 107 499 109
rect 522 123 527 128
rect 522 121 523 123
rect 525 121 527 123
rect 522 119 527 121
rect 475 101 476 103
rect 478 101 479 103
rect 475 99 479 101
rect 442 95 448 96
rect 442 93 445 95
rect 447 93 448 95
rect 442 92 448 93
rect 523 97 527 119
rect 532 128 536 129
rect 532 126 533 128
rect 535 126 536 128
rect 532 120 536 126
rect 532 118 553 120
rect 532 116 537 118
rect 539 116 553 118
rect 532 111 553 112
rect 532 109 533 111
rect 535 109 547 111
rect 549 109 553 111
rect 532 108 553 109
rect 566 130 568 132
rect 564 125 568 130
rect 566 123 568 125
rect 532 104 536 108
rect 564 107 568 123
rect 580 128 584 129
rect 580 126 581 128
rect 583 126 584 128
rect 580 120 584 126
rect 831 136 835 137
rect 822 132 835 136
rect 620 130 625 132
rect 611 128 616 130
rect 580 119 593 120
rect 580 117 585 119
rect 587 117 593 119
rect 580 116 593 117
rect 564 105 565 107
rect 567 105 568 107
rect 564 104 568 105
rect 563 102 568 104
rect 563 100 564 102
rect 566 100 568 102
rect 563 98 568 100
rect 587 111 601 112
rect 587 109 595 111
rect 597 109 601 111
rect 587 108 601 109
rect 611 126 612 128
rect 614 126 616 128
rect 611 121 616 126
rect 611 119 612 121
rect 614 119 616 121
rect 611 117 616 119
rect 587 106 592 108
rect 587 104 589 106
rect 591 104 592 106
rect 587 99 592 104
rect 612 111 616 117
rect 612 109 613 111
rect 615 109 616 111
rect 522 95 529 97
rect 612 97 616 109
rect 522 93 523 95
rect 525 93 526 95
rect 528 93 529 95
rect 522 91 529 93
rect 604 95 612 97
rect 614 95 616 97
rect 604 91 616 95
rect 620 128 622 130
rect 624 128 625 130
rect 620 123 625 128
rect 620 121 622 123
rect 624 121 625 123
rect 620 119 625 121
rect 620 103 624 119
rect 651 119 689 120
rect 651 117 670 119
rect 672 117 689 119
rect 651 116 689 117
rect 651 113 656 116
rect 648 111 656 113
rect 648 109 649 111
rect 651 109 656 111
rect 648 107 656 109
rect 666 111 681 112
rect 666 109 668 111
rect 670 109 672 111
rect 674 109 675 111
rect 677 109 681 111
rect 666 108 681 109
rect 620 101 621 103
rect 623 101 624 103
rect 620 97 624 101
rect 620 95 625 97
rect 668 99 672 108
rect 699 127 705 129
rect 699 125 700 127
rect 702 125 705 127
rect 699 120 705 125
rect 699 118 700 120
rect 702 118 705 120
rect 699 116 705 118
rect 701 111 705 116
rect 701 109 702 111
rect 704 109 705 111
rect 701 96 705 109
rect 620 93 622 95
rect 624 93 625 95
rect 620 91 625 93
rect 699 95 705 96
rect 699 93 700 95
rect 702 93 705 95
rect 699 92 705 93
rect 709 127 715 129
rect 789 130 794 132
rect 789 128 790 130
rect 792 128 794 130
rect 709 125 712 127
rect 714 125 715 127
rect 709 124 715 125
rect 709 122 712 124
rect 714 122 715 124
rect 709 120 715 122
rect 709 118 712 120
rect 714 118 715 120
rect 709 116 715 118
rect 709 96 713 116
rect 725 119 763 120
rect 725 117 760 119
rect 762 117 763 119
rect 725 116 763 117
rect 758 113 763 116
rect 733 111 748 112
rect 733 109 737 111
rect 739 109 744 111
rect 746 109 748 111
rect 733 108 748 109
rect 758 111 766 113
rect 758 109 763 111
rect 765 109 766 111
rect 742 103 746 108
rect 758 107 766 109
rect 789 123 794 128
rect 789 121 790 123
rect 792 121 794 123
rect 789 119 794 121
rect 742 101 743 103
rect 745 101 746 103
rect 742 99 746 101
rect 709 95 715 96
rect 709 93 712 95
rect 714 93 715 95
rect 709 92 715 93
rect 790 97 794 119
rect 799 128 803 129
rect 799 126 800 128
rect 802 126 803 128
rect 799 120 803 126
rect 799 118 820 120
rect 799 116 804 118
rect 806 116 820 118
rect 799 111 820 112
rect 799 109 800 111
rect 802 109 814 111
rect 816 109 820 111
rect 799 108 820 109
rect 833 130 835 132
rect 831 125 835 130
rect 833 123 835 125
rect 799 104 803 108
rect 831 107 835 123
rect 831 105 832 107
rect 834 105 835 107
rect 831 104 835 105
rect 830 102 835 104
rect 830 100 831 102
rect 833 100 835 102
rect 830 98 835 100
rect 789 95 796 97
rect 789 93 790 95
rect 792 93 793 95
rect 795 93 796 95
rect 789 91 796 93
rect 2 85 838 86
rect 2 83 27 85
rect 29 83 37 85
rect 39 83 67 85
rect 69 83 77 85
rect 79 83 296 85
rect 298 83 334 85
rect 336 83 344 85
rect 346 83 563 85
rect 565 83 601 85
rect 603 83 611 85
rect 613 83 830 85
rect 832 83 838 85
rect 2 79 838 83
rect 2 77 763 79
rect 765 77 838 79
rect 2 76 838 77
rect 2 74 131 76
rect 133 74 838 76
rect 2 73 838 74
rect 2 71 27 73
rect 29 71 37 73
rect 39 71 67 73
rect 69 71 77 73
rect 79 71 296 73
rect 298 71 334 73
rect 336 71 344 73
rect 346 71 563 73
rect 565 71 601 73
rect 603 71 611 73
rect 613 71 830 73
rect 832 71 838 73
rect 2 70 838 71
rect 13 55 18 57
rect 13 53 14 55
rect 16 53 18 55
rect 13 48 18 53
rect 30 61 42 65
rect 30 59 38 61
rect 40 59 42 61
rect 13 47 27 48
rect 13 45 21 47
rect 23 45 27 47
rect 13 44 27 45
rect 6 39 19 40
rect 6 37 11 39
rect 13 37 19 39
rect 6 36 19 37
rect 6 35 10 36
rect 6 33 7 35
rect 9 33 10 35
rect 38 42 42 59
rect 53 56 58 57
rect 53 54 55 56
rect 57 54 58 56
rect 53 48 58 54
rect 70 61 82 65
rect 70 59 78 61
rect 80 59 82 61
rect 53 47 67 48
rect 53 45 61 47
rect 63 45 67 47
rect 53 44 67 45
rect 38 40 39 42
rect 41 40 42 42
rect 38 39 42 40
rect 6 27 10 33
rect 37 37 42 39
rect 37 35 38 37
rect 40 35 42 37
rect 37 30 42 35
rect 46 39 59 40
rect 46 38 51 39
rect 46 36 47 38
rect 49 37 51 38
rect 53 37 59 39
rect 49 36 59 37
rect 46 31 50 36
rect 78 47 82 59
rect 78 45 79 47
rect 81 45 82 47
rect 78 39 82 45
rect 37 28 38 30
rect 40 28 42 30
rect 37 26 42 28
rect 77 37 82 39
rect 77 35 78 37
rect 80 35 82 37
rect 77 30 82 35
rect 77 28 78 30
rect 80 28 82 30
rect 77 26 82 28
rect 86 63 91 65
rect 86 61 88 63
rect 90 61 91 63
rect 86 59 91 61
rect 86 55 90 59
rect 86 53 87 55
rect 89 53 90 55
rect 86 37 90 53
rect 165 63 171 64
rect 165 61 166 63
rect 168 61 171 63
rect 165 60 171 61
rect 86 35 91 37
rect 86 33 88 35
rect 90 33 91 35
rect 86 28 91 33
rect 114 47 122 49
rect 134 48 138 57
rect 114 45 115 47
rect 117 45 122 47
rect 114 43 122 45
rect 132 47 147 48
rect 132 45 134 47
rect 136 45 137 47
rect 139 45 141 47
rect 143 45 147 47
rect 132 44 147 45
rect 117 40 122 43
rect 167 47 171 60
rect 167 45 168 47
rect 170 45 171 47
rect 117 39 155 40
rect 117 37 131 39
rect 133 37 155 39
rect 117 36 155 37
rect 167 40 171 45
rect 165 38 171 40
rect 165 36 166 38
rect 168 36 171 38
rect 165 31 171 36
rect 165 29 166 31
rect 168 29 171 31
rect 86 26 88 28
rect 90 26 91 28
rect 86 24 91 26
rect 165 27 171 29
rect 175 63 181 64
rect 175 61 178 63
rect 180 61 181 63
rect 175 60 181 61
rect 255 63 262 65
rect 255 61 256 63
rect 258 61 259 63
rect 261 61 262 63
rect 175 40 179 60
rect 208 55 212 57
rect 208 53 209 55
rect 211 53 212 55
rect 175 38 181 40
rect 175 36 178 38
rect 180 36 181 38
rect 175 34 181 36
rect 175 32 178 34
rect 180 32 181 34
rect 175 31 181 32
rect 175 29 178 31
rect 180 29 181 31
rect 175 27 181 29
rect 208 48 212 53
rect 255 59 262 61
rect 199 47 214 48
rect 199 45 203 47
rect 205 45 210 47
rect 212 45 214 47
rect 199 44 214 45
rect 224 47 232 49
rect 224 45 229 47
rect 231 45 232 47
rect 224 43 232 45
rect 224 42 229 43
rect 224 40 226 42
rect 228 40 229 42
rect 191 36 229 40
rect 256 37 260 59
rect 265 53 269 54
rect 265 51 266 53
rect 268 51 269 53
rect 265 48 269 51
rect 265 47 286 48
rect 265 45 280 47
rect 282 45 286 47
rect 265 44 286 45
rect 296 56 301 58
rect 296 54 297 56
rect 299 54 301 56
rect 296 52 301 54
rect 337 61 349 65
rect 337 59 345 61
rect 347 59 349 61
rect 255 35 260 37
rect 255 33 256 35
rect 258 33 260 35
rect 255 28 260 33
rect 255 26 256 28
rect 258 26 260 28
rect 265 38 270 40
rect 272 38 286 40
rect 265 36 286 38
rect 265 34 269 36
rect 265 32 266 34
rect 268 32 269 34
rect 265 27 269 32
rect 255 24 260 26
rect 297 33 301 52
rect 320 52 325 53
rect 320 50 322 52
rect 324 50 325 52
rect 320 48 325 50
rect 320 47 334 48
rect 320 45 328 47
rect 330 45 334 47
rect 320 44 334 45
rect 299 31 301 33
rect 297 26 301 31
rect 313 39 326 40
rect 313 37 318 39
rect 320 37 326 39
rect 313 36 326 37
rect 313 34 317 36
rect 313 32 314 34
rect 316 32 317 34
rect 345 47 349 59
rect 345 45 346 47
rect 348 45 349 47
rect 345 39 349 45
rect 313 27 317 32
rect 344 37 349 39
rect 344 35 345 37
rect 347 35 349 37
rect 344 30 349 35
rect 299 24 301 26
rect 288 23 301 24
rect 288 21 298 23
rect 300 21 301 23
rect 288 20 301 21
rect 297 19 301 20
rect 344 28 345 30
rect 347 28 349 30
rect 344 26 349 28
rect 353 63 358 65
rect 353 61 355 63
rect 357 61 358 63
rect 353 59 358 61
rect 353 55 357 59
rect 353 53 354 55
rect 356 53 357 55
rect 353 37 357 53
rect 432 63 438 64
rect 432 61 433 63
rect 435 61 438 63
rect 432 60 438 61
rect 353 35 358 37
rect 353 33 355 35
rect 357 33 358 35
rect 353 28 358 33
rect 381 47 389 49
rect 401 48 405 57
rect 381 45 382 47
rect 384 45 389 47
rect 381 43 389 45
rect 399 47 414 48
rect 399 45 401 47
rect 403 45 404 47
rect 406 45 408 47
rect 410 45 414 47
rect 399 44 414 45
rect 384 40 389 43
rect 434 47 438 60
rect 434 45 435 47
rect 437 45 438 47
rect 384 39 422 40
rect 384 37 398 39
rect 400 37 422 39
rect 384 36 422 37
rect 434 40 438 45
rect 432 38 438 40
rect 432 36 433 38
rect 435 36 438 38
rect 432 31 438 36
rect 432 29 433 31
rect 435 29 438 31
rect 353 26 355 28
rect 357 26 358 28
rect 353 24 358 26
rect 432 27 438 29
rect 442 63 448 64
rect 442 61 445 63
rect 447 61 448 63
rect 442 60 448 61
rect 522 63 529 65
rect 522 61 523 63
rect 525 61 526 63
rect 528 61 529 63
rect 442 40 446 60
rect 475 55 479 57
rect 475 53 476 55
rect 478 53 479 55
rect 442 38 448 40
rect 442 36 445 38
rect 447 36 448 38
rect 442 34 448 36
rect 442 32 445 34
rect 447 32 448 34
rect 442 31 448 32
rect 442 29 445 31
rect 447 29 448 31
rect 442 27 448 29
rect 475 48 479 53
rect 522 59 529 61
rect 466 47 481 48
rect 466 45 470 47
rect 472 45 477 47
rect 479 45 481 47
rect 466 44 481 45
rect 491 47 499 49
rect 491 45 496 47
rect 498 45 499 47
rect 491 43 499 45
rect 491 42 496 43
rect 491 40 493 42
rect 495 40 496 42
rect 458 36 496 40
rect 523 37 527 59
rect 532 53 536 54
rect 532 51 533 53
rect 535 51 536 53
rect 532 48 536 51
rect 532 47 553 48
rect 532 45 547 47
rect 549 45 553 47
rect 532 44 553 45
rect 563 56 568 58
rect 563 54 564 56
rect 566 54 568 56
rect 604 61 616 65
rect 604 59 612 61
rect 614 59 616 61
rect 563 52 568 54
rect 522 35 527 37
rect 522 33 523 35
rect 525 33 527 35
rect 522 28 527 33
rect 522 26 523 28
rect 525 26 527 28
rect 532 38 537 40
rect 539 38 553 40
rect 532 36 553 38
rect 532 34 536 36
rect 532 32 533 34
rect 535 32 536 34
rect 532 27 536 32
rect 522 24 527 26
rect 564 33 568 52
rect 587 53 592 54
rect 587 51 589 53
rect 591 51 592 53
rect 587 48 592 51
rect 587 47 601 48
rect 587 45 595 47
rect 597 45 601 47
rect 587 44 601 45
rect 566 31 568 33
rect 564 26 568 31
rect 580 39 593 40
rect 580 37 585 39
rect 587 37 593 39
rect 580 36 593 37
rect 580 34 584 36
rect 580 32 581 34
rect 583 32 584 34
rect 612 47 616 59
rect 612 45 613 47
rect 615 45 616 47
rect 612 39 616 45
rect 580 27 584 32
rect 611 37 616 39
rect 611 35 612 37
rect 614 35 616 37
rect 611 30 616 35
rect 566 24 568 26
rect 555 22 568 24
rect 555 20 565 22
rect 567 20 568 22
rect 564 19 568 20
rect 611 28 612 30
rect 614 28 616 30
rect 611 26 616 28
rect 620 63 625 65
rect 620 61 622 63
rect 624 61 625 63
rect 620 59 625 61
rect 620 55 624 59
rect 620 53 621 55
rect 623 53 624 55
rect 620 37 624 53
rect 699 63 705 64
rect 699 61 700 63
rect 702 61 705 63
rect 699 60 705 61
rect 620 35 625 37
rect 620 33 622 35
rect 624 33 625 35
rect 620 28 625 33
rect 648 47 656 49
rect 668 48 672 57
rect 648 45 649 47
rect 651 45 656 47
rect 648 43 656 45
rect 666 47 681 48
rect 666 45 668 47
rect 670 45 671 47
rect 673 45 675 47
rect 677 45 681 47
rect 666 44 681 45
rect 651 40 656 43
rect 701 47 705 60
rect 701 45 702 47
rect 704 45 705 47
rect 651 39 689 40
rect 651 37 665 39
rect 667 37 689 39
rect 651 36 689 37
rect 701 40 705 45
rect 699 38 705 40
rect 699 36 700 38
rect 702 36 705 38
rect 699 31 705 36
rect 699 29 700 31
rect 702 29 705 31
rect 620 26 622 28
rect 624 26 625 28
rect 620 24 625 26
rect 699 27 705 29
rect 709 63 715 64
rect 709 61 712 63
rect 714 61 715 63
rect 709 60 715 61
rect 789 63 796 65
rect 789 61 790 63
rect 792 61 793 63
rect 795 61 796 63
rect 709 40 713 60
rect 742 55 746 57
rect 742 53 743 55
rect 745 53 746 55
rect 709 38 715 40
rect 709 36 712 38
rect 714 36 715 38
rect 709 34 715 36
rect 709 32 712 34
rect 714 32 715 34
rect 709 31 715 32
rect 709 29 712 31
rect 714 29 715 31
rect 709 27 715 29
rect 742 48 746 53
rect 789 59 796 61
rect 733 47 748 48
rect 733 45 737 47
rect 739 45 744 47
rect 746 45 748 47
rect 733 44 748 45
rect 758 47 766 49
rect 758 45 763 47
rect 765 45 766 47
rect 758 43 766 45
rect 758 42 763 43
rect 758 40 760 42
rect 762 40 763 42
rect 725 36 763 40
rect 790 37 794 59
rect 799 53 803 54
rect 799 51 800 53
rect 802 51 803 53
rect 799 48 803 51
rect 799 47 820 48
rect 799 45 814 47
rect 816 45 820 47
rect 799 44 820 45
rect 830 56 835 58
rect 830 54 831 56
rect 833 54 835 56
rect 830 52 835 54
rect 789 35 794 37
rect 789 33 790 35
rect 792 33 794 35
rect 789 28 794 33
rect 789 26 790 28
rect 792 26 794 28
rect 799 38 804 40
rect 806 38 820 40
rect 799 36 820 38
rect 799 34 803 36
rect 799 32 800 34
rect 802 32 803 34
rect 799 27 803 32
rect 789 24 794 26
rect 831 33 835 52
rect 833 31 835 33
rect 831 26 835 31
rect 833 24 835 26
rect 822 23 835 24
rect 822 21 824 23
rect 826 21 835 23
rect 822 20 835 21
rect 831 19 835 20
rect 2 13 838 14
rect 2 11 37 13
rect 39 11 77 13
rect 79 11 296 13
rect 298 11 344 13
rect 346 11 563 13
rect 565 11 611 13
rect 613 11 830 13
rect 832 11 838 13
rect 2 8 838 11
rect 2 6 25 8
rect 27 6 838 8
rect 2 5 838 6
rect 2 3 832 5
rect 834 3 838 5
rect 2 1 838 3
rect 2 -1 460 1
rect 462 -1 698 1
rect 700 -1 838 1
rect 2 -2 838 -1
rect 424 -8 436 -7
rect 424 -10 432 -8
rect 434 -10 436 -8
rect 424 -13 436 -10
rect 424 -25 429 -13
rect 699 -8 703 -7
rect 690 -9 703 -8
rect 690 -11 700 -9
rect 702 -11 703 -9
rect 690 -12 703 -11
rect 488 -14 493 -12
rect 424 -27 426 -25
rect 428 -27 429 -25
rect 424 -29 429 -27
rect 440 -35 445 -31
rect 440 -37 441 -35
rect 443 -37 445 -35
rect 468 -16 484 -15
rect 468 -18 470 -16
rect 472 -18 484 -16
rect 468 -20 484 -18
rect 480 -25 484 -20
rect 480 -27 481 -25
rect 483 -27 484 -25
rect 440 -38 445 -37
rect 440 -39 442 -38
rect 432 -40 442 -39
rect 444 -40 445 -38
rect 432 -45 445 -40
rect 480 -48 484 -27
rect 460 -49 484 -48
rect 460 -51 462 -49
rect 464 -51 484 -49
rect 460 -52 484 -51
rect 488 -16 490 -14
rect 492 -16 493 -14
rect 488 -21 493 -16
rect 488 -23 490 -21
rect 492 -23 493 -21
rect 488 -25 493 -23
rect 488 -41 492 -25
rect 519 -25 557 -24
rect 519 -27 520 -25
rect 522 -27 557 -25
rect 519 -28 557 -27
rect 519 -31 524 -28
rect 516 -33 524 -31
rect 516 -35 517 -33
rect 519 -35 524 -33
rect 516 -37 524 -35
rect 534 -33 549 -32
rect 534 -35 536 -33
rect 538 -35 540 -33
rect 542 -35 543 -33
rect 545 -35 549 -33
rect 534 -36 549 -35
rect 488 -43 489 -41
rect 491 -43 492 -41
rect 488 -47 492 -43
rect 488 -49 493 -47
rect 536 -45 540 -36
rect 567 -17 573 -15
rect 567 -19 568 -17
rect 570 -19 573 -17
rect 567 -24 573 -19
rect 567 -26 568 -24
rect 570 -26 573 -24
rect 567 -28 573 -26
rect 569 -33 573 -28
rect 569 -35 570 -33
rect 572 -35 573 -33
rect 569 -48 573 -35
rect 488 -51 490 -49
rect 492 -51 493 -49
rect 488 -53 493 -51
rect 567 -49 573 -48
rect 567 -51 568 -49
rect 570 -51 573 -49
rect 567 -52 573 -51
rect 577 -17 583 -15
rect 657 -14 662 -12
rect 657 -16 658 -14
rect 660 -16 662 -14
rect 577 -19 580 -17
rect 582 -19 583 -17
rect 577 -20 583 -19
rect 577 -22 580 -20
rect 582 -22 583 -20
rect 577 -24 583 -22
rect 577 -26 580 -24
rect 582 -26 583 -24
rect 577 -28 583 -26
rect 577 -48 581 -28
rect 593 -28 631 -24
rect 626 -30 628 -28
rect 630 -30 631 -28
rect 626 -31 631 -30
rect 601 -33 616 -32
rect 601 -35 605 -33
rect 607 -35 612 -33
rect 614 -35 616 -33
rect 601 -36 616 -35
rect 626 -33 634 -31
rect 626 -35 631 -33
rect 633 -35 634 -33
rect 610 -41 614 -36
rect 626 -37 634 -35
rect 657 -21 662 -16
rect 657 -23 658 -21
rect 660 -23 662 -21
rect 657 -25 662 -23
rect 610 -43 611 -41
rect 613 -43 614 -41
rect 610 -45 614 -43
rect 577 -49 583 -48
rect 577 -51 580 -49
rect 582 -51 583 -49
rect 577 -52 583 -51
rect 658 -47 662 -25
rect 667 -20 671 -15
rect 667 -22 668 -20
rect 670 -22 671 -20
rect 667 -24 671 -22
rect 667 -26 688 -24
rect 667 -28 672 -26
rect 674 -28 688 -26
rect 667 -33 688 -32
rect 667 -35 682 -33
rect 684 -35 688 -33
rect 667 -36 688 -35
rect 701 -14 703 -12
rect 699 -19 703 -14
rect 701 -21 703 -19
rect 710 -13 715 -7
rect 757 -9 770 -8
rect 757 -11 766 -9
rect 768 -11 770 -9
rect 710 -15 712 -13
rect 714 -15 715 -13
rect 757 -12 770 -11
rect 710 -16 715 -15
rect 710 -17 723 -16
rect 710 -19 720 -17
rect 722 -19 723 -17
rect 710 -20 723 -19
rect 667 -39 671 -36
rect 667 -41 668 -39
rect 670 -41 671 -39
rect 699 -40 703 -21
rect 667 -44 671 -41
rect 698 -42 703 -40
rect 698 -44 699 -42
rect 701 -44 703 -42
rect 698 -46 703 -44
rect 657 -48 662 -47
rect 724 -33 730 -31
rect 724 -35 725 -33
rect 727 -35 730 -33
rect 724 -40 730 -35
rect 717 -41 730 -40
rect 717 -43 719 -41
rect 721 -43 730 -41
rect 742 -25 754 -23
rect 742 -27 747 -25
rect 749 -27 754 -25
rect 742 -28 754 -27
rect 742 -29 752 -28
rect 750 -30 752 -29
rect 750 -37 754 -30
rect 717 -44 730 -43
rect 657 -49 664 -48
rect 657 -51 658 -49
rect 660 -51 661 -49
rect 663 -51 664 -49
rect 766 -45 770 -12
rect 774 -13 779 -7
rect 821 -9 834 -8
rect 821 -11 830 -9
rect 832 -11 834 -9
rect 774 -15 776 -13
rect 778 -15 779 -13
rect 821 -12 834 -11
rect 774 -16 779 -15
rect 774 -17 787 -16
rect 774 -19 776 -17
rect 778 -19 787 -17
rect 774 -20 787 -19
rect 765 -47 770 -45
rect 657 -53 664 -51
rect 765 -49 766 -47
rect 768 -49 770 -47
rect 765 -50 770 -49
rect 765 -51 767 -50
rect 766 -52 767 -51
rect 769 -52 770 -50
rect 788 -33 794 -31
rect 788 -35 789 -33
rect 791 -35 794 -33
rect 788 -36 794 -35
rect 788 -38 790 -36
rect 792 -38 794 -36
rect 788 -40 794 -38
rect 781 -44 794 -40
rect 805 -25 818 -23
rect 805 -27 806 -25
rect 808 -27 818 -25
rect 805 -28 818 -27
rect 805 -29 816 -28
rect 814 -30 816 -29
rect 814 -37 818 -30
rect 830 -17 834 -12
rect 830 -19 831 -17
rect 833 -19 834 -17
rect 830 -45 834 -19
rect 829 -47 834 -45
rect 766 -53 770 -52
rect 829 -49 830 -47
rect 832 -49 834 -47
rect 829 -51 834 -49
rect 830 -53 834 -51
rect 420 -59 838 -58
rect 420 -61 427 -59
rect 429 -61 480 -59
rect 482 -61 698 -59
rect 700 -61 838 -59
rect 420 -65 838 -61
rect 420 -67 762 -65
rect 764 -67 838 -65
rect 420 -71 838 -67
rect 420 -73 427 -71
rect 429 -73 480 -71
rect 482 -73 698 -71
rect 700 -73 838 -71
rect 420 -74 838 -73
rect 460 -81 484 -80
rect 460 -83 462 -81
rect 464 -83 484 -81
rect 460 -84 484 -83
rect 432 -89 445 -87
rect 432 -91 436 -89
rect 438 -91 445 -89
rect 432 -92 445 -91
rect 432 -93 442 -92
rect 440 -94 442 -93
rect 444 -94 445 -92
rect 424 -105 429 -103
rect 424 -107 426 -105
rect 428 -107 429 -105
rect 424 -119 429 -107
rect 440 -101 445 -94
rect 424 -121 425 -119
rect 427 -121 436 -119
rect 424 -125 436 -121
rect 480 -105 484 -84
rect 480 -107 481 -105
rect 483 -107 484 -105
rect 480 -112 484 -107
rect 468 -114 484 -112
rect 468 -116 470 -114
rect 472 -116 484 -114
rect 468 -117 484 -116
rect 488 -81 493 -79
rect 488 -83 490 -81
rect 492 -83 493 -81
rect 488 -85 493 -83
rect 488 -89 492 -85
rect 488 -91 489 -89
rect 491 -91 492 -89
rect 488 -107 492 -91
rect 567 -81 573 -80
rect 567 -83 568 -81
rect 570 -83 573 -81
rect 567 -84 573 -83
rect 488 -109 493 -107
rect 488 -111 490 -109
rect 492 -111 493 -109
rect 488 -116 493 -111
rect 516 -97 524 -95
rect 536 -96 540 -87
rect 516 -99 517 -97
rect 519 -99 524 -97
rect 516 -101 524 -99
rect 534 -97 549 -96
rect 534 -99 536 -97
rect 538 -99 539 -97
rect 541 -99 543 -97
rect 545 -99 549 -97
rect 534 -100 549 -99
rect 519 -104 524 -101
rect 569 -97 573 -84
rect 569 -99 570 -97
rect 572 -99 573 -97
rect 519 -105 557 -104
rect 519 -107 526 -105
rect 528 -107 557 -105
rect 519 -108 557 -107
rect 569 -104 573 -99
rect 567 -106 573 -104
rect 567 -108 568 -106
rect 570 -108 573 -106
rect 567 -113 573 -108
rect 567 -115 568 -113
rect 570 -115 573 -113
rect 488 -118 490 -116
rect 492 -118 493 -116
rect 488 -120 493 -118
rect 567 -117 573 -115
rect 577 -81 583 -80
rect 577 -83 580 -81
rect 582 -83 583 -81
rect 577 -84 583 -83
rect 657 -81 664 -79
rect 657 -83 658 -81
rect 660 -83 661 -81
rect 663 -83 664 -81
rect 577 -104 581 -84
rect 610 -89 614 -87
rect 610 -91 611 -89
rect 613 -91 614 -89
rect 577 -106 583 -104
rect 577 -108 580 -106
rect 582 -108 583 -106
rect 577 -110 583 -108
rect 577 -112 580 -110
rect 582 -112 583 -110
rect 577 -113 583 -112
rect 577 -115 580 -113
rect 582 -115 583 -113
rect 577 -117 583 -115
rect 610 -96 614 -91
rect 657 -84 664 -83
rect 657 -85 662 -84
rect 601 -97 616 -96
rect 601 -99 605 -97
rect 607 -99 612 -97
rect 614 -99 616 -97
rect 601 -100 616 -99
rect 626 -97 634 -95
rect 626 -99 631 -97
rect 633 -99 634 -97
rect 626 -101 634 -99
rect 626 -104 631 -101
rect 593 -105 631 -104
rect 593 -107 628 -105
rect 630 -107 631 -105
rect 593 -108 631 -107
rect 658 -107 662 -85
rect 667 -96 671 -89
rect 667 -97 688 -96
rect 667 -99 668 -97
rect 670 -99 682 -97
rect 684 -99 688 -97
rect 667 -100 688 -99
rect 698 -88 703 -86
rect 698 -90 699 -88
rect 701 -90 703 -88
rect 698 -92 703 -90
rect 657 -109 662 -107
rect 657 -111 658 -109
rect 660 -111 662 -109
rect 657 -116 662 -111
rect 657 -118 658 -116
rect 660 -118 662 -116
rect 667 -106 672 -104
rect 674 -106 688 -104
rect 667 -108 688 -106
rect 667 -114 671 -108
rect 699 -93 703 -92
rect 699 -95 700 -93
rect 702 -95 703 -93
rect 667 -116 668 -114
rect 670 -116 671 -114
rect 667 -117 671 -116
rect 657 -120 662 -118
rect 699 -111 703 -95
rect 766 -81 770 -79
rect 765 -83 770 -81
rect 765 -85 766 -83
rect 768 -85 770 -83
rect 765 -87 770 -85
rect 717 -89 730 -88
rect 717 -91 718 -89
rect 720 -91 730 -89
rect 717 -92 730 -91
rect 724 -97 730 -92
rect 724 -99 725 -97
rect 727 -99 730 -97
rect 724 -101 730 -99
rect 766 -89 770 -87
rect 750 -102 754 -95
rect 766 -91 767 -89
rect 769 -91 770 -89
rect 750 -103 752 -102
rect 743 -104 752 -103
rect 743 -105 754 -104
rect 743 -107 750 -105
rect 752 -107 754 -105
rect 743 -109 754 -107
rect 701 -113 703 -111
rect 699 -118 703 -113
rect 701 -120 703 -118
rect 690 -124 703 -120
rect 699 -125 703 -124
rect 710 -113 723 -112
rect 710 -115 719 -113
rect 721 -115 723 -113
rect 710 -116 723 -115
rect 710 -117 715 -116
rect 710 -119 712 -117
rect 714 -119 715 -117
rect 710 -125 715 -119
rect 766 -120 770 -91
rect 784 -88 790 -85
rect 830 -81 834 -79
rect 829 -83 834 -81
rect 829 -85 830 -83
rect 832 -85 834 -83
rect 829 -87 834 -85
rect 781 -92 794 -88
rect 788 -97 794 -92
rect 788 -99 789 -97
rect 791 -99 794 -97
rect 788 -101 794 -99
rect 814 -102 818 -95
rect 814 -103 816 -102
rect 805 -104 816 -103
rect 805 -105 818 -104
rect 805 -107 806 -105
rect 808 -107 818 -105
rect 805 -109 818 -107
rect 757 -121 770 -120
rect 757 -123 766 -121
rect 768 -123 770 -121
rect 757 -124 770 -123
rect 774 -113 787 -112
rect 774 -115 775 -113
rect 777 -115 787 -113
rect 774 -116 787 -115
rect 774 -117 779 -116
rect 830 -108 834 -87
rect 830 -110 831 -108
rect 833 -110 834 -108
rect 774 -119 776 -117
rect 778 -119 779 -117
rect 774 -125 779 -119
rect 830 -120 834 -110
rect 821 -121 834 -120
rect 821 -123 830 -121
rect 832 -123 834 -121
rect 821 -124 834 -123
rect 420 -131 838 -130
rect 420 -133 460 -131
rect 462 -133 698 -131
rect 700 -133 838 -131
rect 420 -140 838 -133
rect 420 -142 835 -140
rect 837 -142 838 -140
rect 420 -143 838 -142
rect 420 -145 460 -143
rect 462 -145 698 -143
rect 700 -145 838 -143
rect 420 -146 838 -145
rect 424 -157 436 -151
rect 424 -159 429 -157
rect 424 -161 426 -159
rect 428 -161 429 -159
rect 424 -169 429 -161
rect 699 -152 703 -151
rect 690 -156 703 -152
rect 488 -158 493 -156
rect 424 -171 426 -169
rect 428 -171 429 -169
rect 424 -173 429 -171
rect 440 -182 445 -175
rect 468 -160 484 -159
rect 468 -162 470 -160
rect 472 -162 484 -160
rect 468 -164 484 -162
rect 480 -169 484 -164
rect 480 -171 481 -169
rect 483 -171 484 -169
rect 440 -183 442 -182
rect 432 -184 442 -183
rect 444 -184 445 -182
rect 432 -186 445 -184
rect 432 -188 434 -186
rect 436 -188 445 -186
rect 432 -189 445 -188
rect 480 -192 484 -171
rect 460 -193 484 -192
rect 460 -195 462 -193
rect 464 -195 484 -193
rect 460 -196 484 -195
rect 488 -160 490 -158
rect 492 -160 493 -158
rect 488 -165 493 -160
rect 488 -167 490 -165
rect 492 -167 493 -165
rect 488 -169 493 -167
rect 488 -185 492 -169
rect 519 -169 557 -168
rect 519 -171 521 -169
rect 523 -171 557 -169
rect 519 -172 557 -171
rect 519 -175 524 -172
rect 516 -177 524 -175
rect 516 -179 517 -177
rect 519 -179 524 -177
rect 516 -181 524 -179
rect 534 -177 549 -176
rect 534 -179 536 -177
rect 538 -179 540 -177
rect 542 -179 543 -177
rect 545 -179 549 -177
rect 534 -180 549 -179
rect 488 -187 489 -185
rect 491 -187 492 -185
rect 488 -191 492 -187
rect 488 -193 493 -191
rect 536 -189 540 -180
rect 567 -161 573 -159
rect 567 -163 568 -161
rect 570 -163 573 -161
rect 567 -168 573 -163
rect 567 -170 568 -168
rect 570 -170 573 -168
rect 567 -172 573 -170
rect 569 -177 573 -172
rect 569 -179 570 -177
rect 572 -179 573 -177
rect 569 -192 573 -179
rect 488 -195 490 -193
rect 492 -195 493 -193
rect 488 -197 493 -195
rect 567 -193 573 -192
rect 567 -195 568 -193
rect 570 -195 573 -193
rect 567 -196 573 -195
rect 577 -161 583 -159
rect 657 -158 662 -156
rect 657 -160 658 -158
rect 660 -160 662 -158
rect 577 -163 580 -161
rect 582 -163 583 -161
rect 577 -164 583 -163
rect 577 -166 580 -164
rect 582 -166 583 -164
rect 577 -168 583 -166
rect 577 -170 580 -168
rect 582 -170 583 -168
rect 577 -172 583 -170
rect 577 -192 581 -172
rect 593 -172 631 -168
rect 626 -174 628 -172
rect 630 -174 631 -172
rect 626 -175 631 -174
rect 601 -177 616 -176
rect 601 -179 605 -177
rect 607 -179 612 -177
rect 614 -179 616 -177
rect 601 -180 616 -179
rect 626 -177 634 -175
rect 626 -179 631 -177
rect 633 -179 634 -177
rect 610 -185 614 -180
rect 626 -181 634 -179
rect 657 -165 662 -160
rect 657 -167 658 -165
rect 660 -167 662 -165
rect 657 -169 662 -167
rect 610 -187 611 -185
rect 613 -187 614 -185
rect 610 -189 614 -187
rect 577 -193 583 -192
rect 577 -195 580 -193
rect 582 -195 583 -193
rect 577 -196 583 -195
rect 658 -191 662 -169
rect 667 -164 671 -159
rect 667 -166 668 -164
rect 670 -166 671 -164
rect 667 -168 671 -166
rect 667 -170 688 -168
rect 667 -172 672 -170
rect 674 -172 688 -170
rect 667 -177 688 -176
rect 667 -179 682 -177
rect 684 -179 688 -177
rect 667 -180 688 -179
rect 701 -158 703 -156
rect 699 -163 703 -158
rect 701 -165 703 -163
rect 710 -157 715 -151
rect 757 -153 770 -152
rect 757 -155 766 -153
rect 768 -155 770 -153
rect 710 -159 712 -157
rect 714 -159 715 -157
rect 757 -156 770 -155
rect 710 -160 715 -159
rect 710 -161 723 -160
rect 710 -163 718 -161
rect 720 -163 723 -161
rect 710 -164 723 -163
rect 667 -183 671 -180
rect 667 -185 668 -183
rect 670 -185 671 -183
rect 699 -182 703 -165
rect 699 -184 700 -182
rect 702 -184 703 -182
rect 667 -187 671 -185
rect 698 -186 703 -184
rect 698 -188 699 -186
rect 701 -188 703 -186
rect 698 -190 703 -188
rect 724 -177 730 -175
rect 724 -179 725 -177
rect 727 -179 730 -177
rect 724 -184 730 -179
rect 717 -185 730 -184
rect 717 -187 718 -185
rect 720 -187 730 -185
rect 742 -169 754 -167
rect 742 -171 745 -169
rect 747 -171 754 -169
rect 742 -172 754 -171
rect 742 -173 752 -172
rect 750 -174 752 -173
rect 750 -181 754 -174
rect 766 -169 770 -156
rect 774 -157 779 -151
rect 821 -153 834 -152
rect 821 -155 830 -153
rect 832 -155 834 -153
rect 774 -159 776 -157
rect 778 -159 779 -157
rect 821 -156 834 -155
rect 774 -160 779 -159
rect 774 -161 787 -160
rect 774 -163 776 -161
rect 778 -163 787 -161
rect 774 -164 787 -163
rect 766 -171 767 -169
rect 769 -171 770 -169
rect 717 -188 730 -187
rect 657 -193 664 -191
rect 657 -195 658 -193
rect 660 -195 661 -193
rect 663 -195 664 -193
rect 766 -189 770 -171
rect 765 -191 770 -189
rect 657 -197 664 -195
rect 765 -193 766 -191
rect 768 -193 770 -191
rect 765 -195 770 -193
rect 788 -177 794 -175
rect 788 -179 789 -177
rect 791 -179 794 -177
rect 788 -184 794 -179
rect 781 -188 794 -184
rect 806 -170 818 -167
rect 806 -172 807 -170
rect 809 -172 818 -170
rect 806 -173 816 -172
rect 814 -174 816 -173
rect 814 -181 818 -174
rect 830 -168 834 -156
rect 830 -170 831 -168
rect 833 -170 834 -168
rect 784 -191 790 -188
rect 830 -189 834 -170
rect 829 -191 834 -189
rect 766 -197 770 -195
rect 829 -193 830 -191
rect 832 -193 834 -191
rect 829 -195 834 -193
rect 830 -197 834 -195
rect 420 -203 838 -202
rect 420 -205 427 -203
rect 429 -205 480 -203
rect 482 -205 698 -203
rect 700 -205 838 -203
rect 420 -209 838 -205
rect 420 -211 765 -209
rect 767 -211 838 -209
rect 420 -215 838 -211
rect 420 -217 427 -215
rect 429 -217 480 -215
rect 482 -217 698 -215
rect 700 -217 838 -215
rect 420 -218 838 -217
rect 460 -225 484 -224
rect 460 -227 462 -225
rect 464 -227 484 -225
rect 460 -228 484 -227
rect 432 -232 445 -231
rect 432 -234 435 -232
rect 437 -234 445 -232
rect 432 -236 445 -234
rect 432 -237 442 -236
rect 440 -238 442 -237
rect 444 -238 445 -236
rect 424 -249 429 -247
rect 424 -251 426 -249
rect 428 -251 429 -249
rect 424 -255 429 -251
rect 440 -245 445 -238
rect 424 -257 426 -255
rect 428 -257 429 -255
rect 424 -263 429 -257
rect 424 -269 436 -263
rect 480 -249 484 -228
rect 480 -251 481 -249
rect 483 -251 484 -249
rect 480 -256 484 -251
rect 468 -258 484 -256
rect 468 -260 470 -258
rect 472 -260 484 -258
rect 468 -261 484 -260
rect 488 -225 493 -223
rect 488 -227 490 -225
rect 492 -227 493 -225
rect 488 -229 493 -227
rect 488 -233 492 -229
rect 488 -235 489 -233
rect 491 -235 492 -233
rect 488 -251 492 -235
rect 567 -225 573 -224
rect 567 -227 568 -225
rect 570 -227 573 -225
rect 567 -228 573 -227
rect 488 -253 493 -251
rect 488 -255 490 -253
rect 492 -255 493 -253
rect 488 -260 493 -255
rect 516 -241 524 -239
rect 536 -240 540 -231
rect 516 -243 517 -241
rect 519 -243 524 -241
rect 516 -245 524 -243
rect 534 -241 549 -240
rect 534 -243 536 -241
rect 538 -243 540 -241
rect 542 -243 543 -241
rect 545 -243 549 -241
rect 534 -244 549 -243
rect 519 -248 524 -245
rect 569 -241 573 -228
rect 569 -243 570 -241
rect 572 -243 573 -241
rect 519 -249 557 -248
rect 519 -251 531 -249
rect 533 -251 557 -249
rect 519 -252 557 -251
rect 569 -248 573 -243
rect 567 -250 573 -248
rect 567 -252 568 -250
rect 570 -252 573 -250
rect 567 -257 573 -252
rect 567 -259 568 -257
rect 570 -259 573 -257
rect 488 -262 490 -260
rect 492 -262 493 -260
rect 488 -264 493 -262
rect 567 -261 573 -259
rect 577 -225 583 -224
rect 577 -227 580 -225
rect 582 -227 583 -225
rect 577 -228 583 -227
rect 657 -225 664 -223
rect 657 -227 658 -225
rect 660 -227 661 -225
rect 663 -227 664 -225
rect 577 -248 581 -228
rect 610 -233 614 -231
rect 610 -235 611 -233
rect 613 -235 614 -233
rect 577 -250 583 -248
rect 577 -252 580 -250
rect 582 -252 583 -250
rect 577 -254 583 -252
rect 577 -256 580 -254
rect 582 -256 583 -254
rect 577 -257 583 -256
rect 577 -259 580 -257
rect 582 -259 583 -257
rect 577 -261 583 -259
rect 610 -240 614 -235
rect 657 -229 664 -227
rect 601 -241 616 -240
rect 601 -243 605 -241
rect 607 -243 612 -241
rect 614 -243 616 -241
rect 601 -244 616 -243
rect 626 -241 634 -239
rect 626 -243 631 -241
rect 633 -243 634 -241
rect 626 -245 634 -243
rect 626 -248 631 -245
rect 593 -249 631 -248
rect 593 -251 622 -249
rect 624 -251 631 -249
rect 593 -252 631 -251
rect 658 -251 662 -229
rect 667 -240 671 -233
rect 667 -241 688 -240
rect 667 -243 668 -241
rect 670 -243 682 -241
rect 684 -243 688 -241
rect 667 -244 688 -243
rect 698 -232 703 -230
rect 698 -234 699 -232
rect 701 -234 703 -232
rect 698 -236 703 -234
rect 657 -253 662 -251
rect 657 -255 658 -253
rect 660 -255 662 -253
rect 657 -260 662 -255
rect 657 -262 658 -260
rect 660 -262 662 -260
rect 667 -250 672 -248
rect 674 -250 688 -248
rect 667 -252 688 -250
rect 667 -254 671 -252
rect 667 -256 668 -254
rect 670 -256 671 -254
rect 699 -237 703 -236
rect 699 -239 700 -237
rect 702 -239 703 -237
rect 667 -261 671 -256
rect 657 -264 662 -262
rect 699 -255 703 -239
rect 766 -225 770 -223
rect 765 -227 770 -225
rect 765 -229 766 -227
rect 768 -229 770 -227
rect 765 -231 770 -229
rect 717 -233 730 -232
rect 717 -235 718 -233
rect 720 -235 730 -233
rect 717 -236 730 -235
rect 724 -241 730 -236
rect 724 -243 725 -241
rect 727 -243 730 -241
rect 724 -245 730 -243
rect 750 -246 754 -239
rect 750 -247 752 -246
rect 742 -248 752 -247
rect 742 -249 754 -248
rect 742 -251 749 -249
rect 751 -251 754 -249
rect 742 -253 754 -251
rect 701 -257 703 -255
rect 699 -262 703 -257
rect 701 -264 703 -262
rect 690 -268 703 -264
rect 699 -269 703 -268
rect 710 -260 723 -256
rect 710 -261 715 -260
rect 766 -253 770 -231
rect 784 -232 790 -229
rect 830 -225 834 -223
rect 829 -227 834 -225
rect 829 -229 830 -227
rect 832 -229 834 -227
rect 829 -231 834 -229
rect 781 -236 794 -232
rect 788 -241 794 -236
rect 788 -243 789 -241
rect 791 -243 794 -241
rect 788 -245 794 -243
rect 814 -246 818 -239
rect 814 -247 816 -246
rect 806 -248 816 -247
rect 806 -249 818 -248
rect 806 -251 814 -249
rect 816 -251 818 -249
rect 806 -253 818 -251
rect 766 -255 767 -253
rect 769 -255 770 -253
rect 710 -263 712 -261
rect 714 -263 715 -261
rect 710 -266 715 -263
rect 766 -264 770 -255
rect 757 -265 770 -264
rect 710 -268 712 -266
rect 714 -268 715 -266
rect 757 -267 766 -265
rect 768 -267 770 -265
rect 757 -268 770 -267
rect 774 -260 787 -256
rect 774 -261 779 -260
rect 830 -249 834 -231
rect 830 -251 831 -249
rect 833 -251 834 -249
rect 774 -263 776 -261
rect 778 -263 779 -261
rect 774 -266 779 -263
rect 830 -264 834 -251
rect 821 -265 834 -264
rect 774 -268 776 -266
rect 778 -268 779 -266
rect 821 -267 830 -265
rect 832 -267 834 -265
rect 821 -268 834 -267
rect 710 -269 715 -268
rect 774 -269 779 -268
rect 420 -275 838 -274
rect 420 -277 460 -275
rect 462 -277 698 -275
rect 700 -277 838 -275
rect 420 -279 838 -277
rect 420 -280 529 -279
rect 420 -282 461 -280
rect 463 -281 529 -280
rect 531 -281 612 -279
rect 614 -281 709 -279
rect 711 -281 773 -279
rect 775 -281 838 -279
rect 463 -282 838 -281
rect 460 -283 469 -282
<< alu2 >>
rect 25 294 34 295
rect 25 293 31 294
rect 25 291 26 293
rect 28 292 31 293
rect 33 292 34 294
rect 28 291 34 292
rect 25 290 34 291
rect 158 294 167 295
rect 158 293 164 294
rect 158 291 159 293
rect 161 292 164 293
rect 166 292 167 294
rect 161 291 167 292
rect 158 290 167 291
rect 398 294 407 295
rect 398 293 404 294
rect 398 291 399 293
rect 401 292 404 293
rect 406 292 407 294
rect 401 291 407 292
rect 398 290 407 291
rect 583 294 592 295
rect 583 293 589 294
rect 583 291 584 293
rect 586 292 589 293
rect 591 292 592 294
rect 586 291 592 292
rect 583 290 592 291
rect 775 294 784 295
rect 775 293 781 294
rect 775 291 776 293
rect 778 292 781 293
rect 783 292 784 294
rect 778 291 784 292
rect 775 290 784 291
rect 46 272 56 273
rect 46 270 47 272
rect 49 270 53 272
rect 55 270 56 272
rect 46 269 56 270
rect 181 272 269 273
rect 181 270 266 272
rect 268 270 269 272
rect 181 269 269 270
rect 304 272 317 273
rect 304 270 305 272
rect 307 270 314 272
rect 316 270 317 272
rect 304 269 317 270
rect 448 272 536 273
rect 448 270 533 272
rect 535 270 536 272
rect 448 269 536 270
rect 573 272 584 273
rect 573 270 574 272
rect 576 270 581 272
rect 583 270 584 272
rect 573 269 584 270
rect 715 272 803 273
rect 715 270 800 272
rect 802 270 803 272
rect 715 269 803 270
rect 177 268 185 269
rect 0 266 10 267
rect 0 264 1 266
rect 3 264 7 266
rect 9 264 10 266
rect 177 266 178 268
rect 180 266 185 268
rect 177 265 185 266
rect 444 268 452 269
rect 444 266 445 268
rect 447 266 452 268
rect 444 265 452 266
rect 711 268 719 269
rect 711 266 712 268
rect 714 266 719 268
rect 711 265 719 266
rect 0 263 10 264
rect 43 263 122 264
rect 43 261 119 263
rect 121 261 122 263
rect 38 260 122 261
rect 207 263 215 264
rect 207 261 208 263
rect 210 261 211 263
rect 213 261 215 263
rect 207 260 215 261
rect 332 263 389 264
rect 332 261 333 263
rect 335 261 386 263
rect 388 261 389 263
rect 332 260 389 261
rect 474 263 482 264
rect 474 261 475 263
rect 477 261 478 263
rect 480 261 482 263
rect 474 260 482 261
rect 599 263 656 264
rect 599 261 600 263
rect 602 261 653 263
rect 655 261 656 263
rect 599 260 656 261
rect 741 263 749 264
rect 741 261 742 263
rect 744 261 745 263
rect 747 261 749 263
rect 741 260 749 261
rect 38 258 39 260
rect 41 258 47 260
rect 38 257 47 258
rect 78 255 140 256
rect 78 253 79 255
rect 81 253 137 255
rect 139 253 140 255
rect 78 252 140 253
rect 167 255 270 256
rect 167 253 168 255
rect 170 253 266 255
rect 268 253 270 255
rect 167 252 270 253
rect 345 255 407 256
rect 345 253 346 255
rect 348 253 404 255
rect 406 253 407 255
rect 345 252 407 253
rect 434 255 537 256
rect 434 253 435 255
rect 437 253 533 255
rect 535 253 537 255
rect 434 252 537 253
rect 612 255 674 256
rect 612 253 613 255
rect 615 253 671 255
rect 673 253 674 255
rect 612 252 674 253
rect 701 255 804 256
rect 701 253 702 255
rect 704 253 800 255
rect 802 253 804 255
rect 701 252 804 253
rect 297 251 305 252
rect 42 249 58 250
rect 42 247 43 249
rect 45 247 55 249
rect 57 247 58 249
rect 297 249 298 251
rect 300 249 302 251
rect 304 249 305 251
rect 564 251 572 252
rect 297 248 305 249
rect 309 249 325 250
rect 13 246 24 247
rect 13 244 15 246
rect 17 244 21 246
rect 23 244 24 246
rect 42 245 58 247
rect 86 247 212 248
rect 86 245 87 247
rect 89 245 209 247
rect 211 245 212 247
rect 309 247 310 249
rect 312 247 322 249
rect 324 247 325 249
rect 564 249 565 251
rect 567 249 569 251
rect 571 249 572 251
rect 831 251 839 252
rect 564 248 572 249
rect 576 249 592 250
rect 309 245 325 247
rect 353 247 479 248
rect 353 245 354 247
rect 356 245 476 247
rect 478 245 479 247
rect 576 247 577 249
rect 579 247 589 249
rect 591 247 592 249
rect 831 249 832 251
rect 834 249 836 251
rect 838 249 839 251
rect 831 248 839 249
rect 86 244 212 245
rect 256 244 265 245
rect 353 244 479 245
rect 523 245 532 246
rect 576 245 592 247
rect 620 247 746 248
rect 620 245 621 247
rect 623 245 743 247
rect 745 245 746 247
rect 13 243 24 244
rect 256 242 257 244
rect 259 242 262 244
rect 264 242 265 244
rect 523 243 524 245
rect 526 243 529 245
rect 531 243 532 245
rect 620 244 746 245
rect 754 245 794 246
rect 523 242 532 243
rect 754 243 755 245
rect 757 243 791 245
rect 793 243 794 245
rect 754 242 794 243
rect 256 241 265 242
rect 210 226 217 227
rect 210 224 211 226
rect 213 224 214 226
rect 216 224 217 226
rect 210 223 217 224
rect 477 226 484 227
rect 477 224 478 226
rect 480 224 481 226
rect 483 224 484 226
rect 477 223 484 224
rect 744 226 751 227
rect 744 224 745 226
rect 747 224 748 226
rect 750 224 751 226
rect 744 223 751 224
rect 768 223 776 226
rect 768 221 769 223
rect 771 221 773 223
rect 775 221 776 223
rect 768 218 776 221
rect 788 208 796 209
rect 258 207 336 208
rect 258 205 259 207
rect 261 205 333 207
rect 335 205 336 207
rect 258 204 336 205
rect 525 207 603 208
rect 525 205 526 207
rect 528 205 600 207
rect 602 205 603 207
rect 788 206 789 208
rect 791 206 793 208
rect 795 206 796 208
rect 788 205 796 206
rect 525 204 603 205
rect 86 199 212 200
rect 353 199 479 200
rect 53 197 65 198
rect 0 195 18 196
rect 0 193 1 195
rect 3 193 15 195
rect 17 193 18 195
rect 53 195 55 197
rect 57 195 62 197
rect 64 195 65 197
rect 86 197 87 199
rect 89 197 209 199
rect 211 197 212 199
rect 289 198 325 199
rect 86 196 212 197
rect 216 197 269 198
rect 53 194 65 195
rect 216 195 266 197
rect 268 195 269 197
rect 289 196 290 198
rect 292 196 322 198
rect 324 196 325 198
rect 353 197 354 199
rect 356 197 476 199
rect 478 197 479 199
rect 620 199 746 200
rect 353 196 479 197
rect 483 197 536 198
rect 620 197 621 199
rect 623 197 743 199
rect 745 197 746 199
rect 289 195 325 196
rect 483 195 533 197
rect 535 195 536 197
rect 216 194 269 195
rect 483 194 536 195
rect 554 196 591 197
rect 620 196 746 197
rect 750 197 803 198
rect 554 194 555 196
rect 557 194 588 196
rect 590 194 591 196
rect 0 192 18 193
rect 216 192 220 194
rect 483 192 487 194
rect 554 193 591 194
rect 750 195 800 197
rect 802 195 803 197
rect 750 194 803 195
rect 750 192 754 194
rect 78 191 140 192
rect 78 189 79 191
rect 81 189 137 191
rect 139 189 140 191
rect 78 188 140 189
rect 167 191 220 192
rect 167 189 168 191
rect 170 189 220 191
rect 167 188 220 189
rect 345 191 407 192
rect 345 189 346 191
rect 348 189 404 191
rect 406 189 407 191
rect 345 188 407 189
rect 434 191 487 192
rect 434 189 435 191
rect 437 189 487 191
rect 434 188 487 189
rect 612 191 674 192
rect 612 189 613 191
rect 615 189 671 191
rect 673 189 674 191
rect 612 188 674 189
rect 701 191 754 192
rect 701 189 702 191
rect 704 189 754 191
rect 701 188 754 189
rect 225 186 305 187
rect 225 184 226 186
rect 228 184 302 186
rect 304 184 305 186
rect 492 186 572 187
rect 492 184 493 186
rect 495 184 569 186
rect 571 184 572 186
rect 759 186 839 187
rect 759 184 760 186
rect 762 184 836 186
rect 838 184 839 186
rect 38 183 135 184
rect 225 183 305 184
rect 320 183 402 184
rect 492 183 572 184
rect 576 183 669 184
rect 759 183 839 184
rect 38 181 39 183
rect 41 181 132 183
rect 134 181 135 183
rect 38 180 135 181
rect 320 181 321 183
rect 323 181 399 183
rect 401 181 402 183
rect 320 180 402 181
rect 576 181 589 183
rect 591 181 666 183
rect 668 181 669 183
rect 576 180 669 181
rect 177 178 269 179
rect 177 176 178 178
rect 180 176 266 178
rect 268 176 269 178
rect 444 178 536 179
rect 444 176 445 178
rect 447 176 533 178
rect 535 176 536 178
rect 711 178 803 179
rect 711 176 712 178
rect 714 176 800 178
rect 802 176 803 178
rect 42 175 50 176
rect 177 175 269 176
rect 309 175 317 176
rect 444 175 536 176
rect 576 175 584 176
rect 711 175 803 176
rect 6 174 18 175
rect 6 172 7 174
rect 9 172 15 174
rect 17 172 18 174
rect 42 173 43 175
rect 45 173 47 175
rect 49 173 50 175
rect 42 172 50 173
rect 309 173 310 175
rect 312 173 314 175
rect 316 173 317 175
rect 309 172 317 173
rect 576 173 577 175
rect 579 173 581 175
rect 583 173 584 175
rect 576 172 584 173
rect 6 171 18 172
rect 289 167 293 168
rect 289 165 290 167
rect 292 165 293 167
rect 6 145 12 146
rect 6 143 8 145
rect 10 143 12 145
rect 6 142 12 143
rect 7 138 12 142
rect -10 135 12 138
rect -10 133 -9 135
rect -7 133 12 135
rect -10 132 12 133
rect 46 128 67 129
rect 46 126 47 128
rect 49 126 64 128
rect 66 126 67 128
rect 46 125 67 126
rect 217 128 269 129
rect 217 126 266 128
rect 268 126 269 128
rect 217 125 269 126
rect 177 124 221 125
rect 0 122 10 123
rect 0 120 1 122
rect 3 120 7 122
rect 9 120 10 122
rect 177 122 178 124
rect 180 122 221 124
rect 177 121 221 122
rect 289 120 293 165
rect 556 167 560 168
rect 556 165 557 167
rect 559 165 560 167
rect 484 128 536 129
rect 484 126 533 128
rect 535 126 536 128
rect 484 125 536 126
rect 298 124 317 125
rect 298 122 299 124
rect 301 122 314 124
rect 316 122 317 124
rect 298 121 317 122
rect 444 124 488 125
rect 444 122 445 124
rect 447 122 488 124
rect 444 121 488 122
rect 556 120 560 165
rect 823 167 827 168
rect 823 165 824 167
rect 826 165 827 167
rect 567 128 584 129
rect 567 126 568 128
rect 570 126 581 128
rect 583 126 584 128
rect 567 125 584 126
rect 751 128 803 129
rect 751 126 800 128
rect 802 126 803 128
rect 751 125 803 126
rect 711 124 755 125
rect 711 122 712 124
rect 714 122 755 124
rect 711 121 755 122
rect 823 120 827 165
rect 832 154 837 155
rect 832 152 834 154
rect 836 152 837 154
rect 832 149 837 152
rect 832 147 833 149
rect 835 147 837 149
rect 832 146 837 147
rect 0 119 10 120
rect 37 119 139 120
rect 37 117 39 119
rect 41 117 136 119
rect 138 117 139 119
rect 37 116 139 117
rect 225 119 293 120
rect 225 117 226 119
rect 228 117 293 119
rect 225 116 293 117
rect 333 119 406 120
rect 333 117 334 119
rect 336 117 403 119
rect 405 117 406 119
rect 333 116 406 117
rect 492 119 560 120
rect 492 117 493 119
rect 495 117 560 119
rect 492 116 560 117
rect 599 119 673 120
rect 599 117 600 119
rect 602 117 670 119
rect 672 117 673 119
rect 599 116 673 117
rect 759 119 827 120
rect 759 117 760 119
rect 762 117 827 119
rect 759 116 827 117
rect 78 111 141 112
rect 78 109 79 111
rect 81 109 138 111
rect 140 109 141 111
rect 78 108 141 109
rect 167 111 270 112
rect 167 109 168 111
rect 170 109 266 111
rect 268 109 270 111
rect 167 108 270 109
rect 345 111 408 112
rect 345 109 346 111
rect 348 109 405 111
rect 407 109 408 111
rect 345 108 408 109
rect 434 111 537 112
rect 434 109 435 111
rect 437 109 533 111
rect 535 109 537 111
rect 434 108 537 109
rect 612 111 675 112
rect 612 109 613 111
rect 615 109 672 111
rect 674 109 675 111
rect 612 108 675 109
rect 701 111 804 112
rect 701 109 702 111
rect 704 109 800 111
rect 802 109 804 111
rect 701 108 804 109
rect 297 107 305 108
rect 564 107 572 108
rect 831 107 839 108
rect 42 106 58 107
rect 42 104 43 106
rect 45 104 55 106
rect 57 104 58 106
rect 297 105 298 107
rect 300 105 302 107
rect 304 105 305 107
rect 297 104 305 105
rect 309 106 325 107
rect 309 104 310 106
rect 312 104 322 106
rect 324 104 325 106
rect 564 105 565 107
rect 567 105 569 107
rect 571 105 572 107
rect 564 104 572 105
rect 576 106 592 107
rect 576 104 577 106
rect 579 104 589 106
rect 591 104 592 106
rect 831 105 832 107
rect 834 105 836 107
rect 838 105 839 107
rect 831 104 839 105
rect 13 103 26 104
rect 42 103 58 104
rect 86 103 212 104
rect 309 103 325 104
rect 353 103 479 104
rect 576 103 592 104
rect 620 103 746 104
rect 13 101 14 103
rect 16 101 23 103
rect 25 101 26 103
rect 13 100 26 101
rect 86 101 87 103
rect 89 101 209 103
rect 211 101 212 103
rect 86 100 212 101
rect 353 101 354 103
rect 356 101 476 103
rect 478 101 479 103
rect 353 100 479 101
rect 620 101 621 103
rect 623 101 743 103
rect 745 101 746 103
rect 620 100 746 101
rect 258 95 324 96
rect 258 93 259 95
rect 261 93 321 95
rect 323 93 324 95
rect 258 91 324 93
rect 525 95 592 96
rect 525 93 526 95
rect 528 93 589 95
rect 591 93 592 95
rect 525 92 592 93
rect 792 95 804 96
rect 792 93 793 95
rect 795 93 801 95
rect 803 93 804 95
rect 792 92 804 93
rect 762 79 770 82
rect 762 77 763 79
rect 765 77 767 79
rect 769 77 770 79
rect 126 76 134 77
rect 126 74 127 76
rect 129 74 131 76
rect 133 74 134 76
rect 762 74 770 77
rect 126 73 134 74
rect 525 64 604 65
rect 258 63 337 64
rect 258 61 259 63
rect 261 61 334 63
rect 336 61 337 63
rect 258 60 337 61
rect 525 63 601 64
rect 525 61 526 63
rect 528 62 601 63
rect 603 62 604 64
rect 528 61 604 62
rect 525 60 604 61
rect 792 63 815 64
rect 792 61 793 63
rect 795 61 811 63
rect 813 61 815 63
rect 792 60 815 61
rect 54 56 65 57
rect 13 55 34 56
rect 13 53 14 55
rect 16 53 31 55
rect 33 53 34 55
rect 54 54 55 56
rect 57 54 62 56
rect 64 54 65 56
rect 54 53 65 54
rect 86 55 212 56
rect 86 53 87 55
rect 89 53 209 55
rect 211 53 212 55
rect 353 55 479 56
rect 13 52 34 53
rect 86 52 212 53
rect 216 53 269 54
rect 353 53 354 55
rect 356 53 476 55
rect 478 53 479 55
rect 620 55 746 56
rect 216 51 266 53
rect 268 51 269 53
rect 42 50 50 51
rect 42 48 43 50
rect 45 48 50 50
rect 216 50 269 51
rect 289 52 325 53
rect 353 52 479 53
rect 483 53 536 54
rect 289 50 290 52
rect 292 50 322 52
rect 324 50 325 52
rect 216 48 220 50
rect 289 49 325 50
rect 483 51 533 53
rect 535 51 536 53
rect 483 50 536 51
rect 551 53 592 54
rect 551 51 552 53
rect 554 51 589 53
rect 591 51 592 53
rect 620 53 621 55
rect 623 53 743 55
rect 745 53 746 55
rect 620 52 746 53
rect 750 53 803 54
rect 551 50 592 51
rect 750 51 800 53
rect 802 51 803 53
rect 750 50 803 51
rect 483 48 487 50
rect 750 48 754 50
rect 42 47 50 48
rect 38 42 42 43
rect 38 40 39 42
rect 41 40 42 42
rect 0 35 10 36
rect 0 33 1 35
rect 3 33 7 35
rect 9 33 10 35
rect 0 32 10 33
rect 38 22 42 40
rect 46 38 50 47
rect 78 47 140 48
rect 78 45 79 47
rect 81 45 137 47
rect 139 45 140 47
rect 78 44 140 45
rect 167 47 220 48
rect 167 45 168 47
rect 170 45 220 47
rect 167 44 220 45
rect 345 47 407 48
rect 345 45 346 47
rect 348 45 404 47
rect 406 45 407 47
rect 345 44 407 45
rect 434 47 487 48
rect 434 45 435 47
rect 437 45 487 47
rect 434 44 487 45
rect 612 47 674 48
rect 612 45 613 47
rect 615 45 671 47
rect 673 45 674 47
rect 612 44 674 45
rect 701 47 754 48
rect 701 45 702 47
rect 704 45 754 47
rect 701 44 754 45
rect 225 42 305 43
rect 225 40 226 42
rect 228 40 302 42
rect 304 40 305 42
rect 492 42 572 43
rect 492 40 493 42
rect 495 40 569 42
rect 571 40 572 42
rect 759 42 839 43
rect 759 40 760 42
rect 762 40 836 42
rect 838 40 839 42
rect 46 36 47 38
rect 49 36 50 38
rect 126 39 134 40
rect 225 39 305 40
rect 393 39 401 40
rect 492 39 572 40
rect 660 39 668 40
rect 759 39 839 40
rect 126 37 127 39
rect 129 37 131 39
rect 133 37 134 39
rect 126 36 134 37
rect 393 37 394 39
rect 396 37 398 39
rect 400 37 401 39
rect 393 36 401 37
rect 660 37 661 39
rect 663 37 665 39
rect 667 37 668 39
rect 660 36 668 37
rect 46 35 50 36
rect 177 34 269 35
rect 177 32 178 34
rect 180 32 266 34
rect 268 32 269 34
rect 177 31 269 32
rect 309 34 317 35
rect 309 32 310 34
rect 312 32 314 34
rect 316 32 317 34
rect 309 31 317 32
rect 444 34 536 35
rect 444 32 445 34
rect 447 32 533 34
rect 535 32 536 34
rect 444 31 536 32
rect 576 34 584 35
rect 576 32 577 34
rect 579 32 581 34
rect 583 32 584 34
rect 576 31 584 32
rect 711 34 803 35
rect 711 32 712 34
rect 714 32 800 34
rect 802 32 803 34
rect 711 31 803 32
rect 38 20 39 22
rect 41 20 42 22
rect 297 23 397 24
rect 820 23 827 24
rect 297 21 298 23
rect 300 21 394 23
rect 396 21 397 23
rect 297 20 397 21
rect 564 22 664 23
rect 564 20 565 22
rect 567 20 661 22
rect 663 20 664 22
rect 820 21 821 23
rect 823 21 824 23
rect 826 21 827 23
rect 820 20 827 21
rect 38 19 42 20
rect 564 19 664 20
rect 831 10 836 11
rect 19 8 28 9
rect 19 6 20 8
rect 22 6 25 8
rect 27 6 28 8
rect 19 5 28 6
rect 831 8 833 10
rect 835 8 836 10
rect 831 5 836 8
rect 38 4 408 5
rect 38 2 39 4
rect 41 2 405 4
rect 407 2 408 4
rect 831 3 832 5
rect 834 3 836 5
rect 831 2 836 3
rect 38 1 408 2
rect 389 -8 580 -7
rect 389 -10 390 -8
rect 392 -10 432 -8
rect 434 -10 577 -8
rect 579 -10 580 -8
rect 389 -11 580 -10
rect 699 -9 715 -8
rect 699 -11 700 -9
rect 702 -11 715 -9
rect 699 -12 715 -11
rect 579 -20 671 -19
rect 579 -22 580 -20
rect 582 -22 668 -20
rect 670 -22 671 -20
rect 579 -23 671 -22
rect 480 -25 523 -24
rect 480 -27 481 -25
rect 483 -27 520 -25
rect 522 -27 523 -25
rect 480 -28 523 -27
rect 540 -27 544 -26
rect 540 -29 541 -27
rect 543 -29 544 -27
rect 540 -32 544 -29
rect 627 -28 707 -27
rect 627 -30 628 -28
rect 630 -30 704 -28
rect 706 -30 707 -28
rect 627 -31 707 -30
rect 711 -32 715 -12
rect 719 -17 783 -16
rect 719 -19 720 -17
rect 722 -19 730 -17
rect 732 -19 776 -17
rect 778 -19 783 -17
rect 719 -20 783 -19
rect 830 -17 834 -16
rect 830 -19 831 -17
rect 833 -19 834 -17
rect 830 -20 834 -19
rect 830 -22 831 -20
rect 833 -22 834 -20
rect 830 -23 834 -22
rect 745 -25 754 -24
rect 745 -27 747 -25
rect 749 -27 751 -25
rect 753 -27 754 -25
rect 745 -28 754 -27
rect 788 -25 810 -24
rect 788 -26 806 -25
rect 788 -28 789 -26
rect 791 -27 806 -26
rect 808 -27 810 -25
rect 791 -28 810 -27
rect 788 -29 810 -28
rect 539 -33 544 -32
rect 417 -35 444 -34
rect 417 -37 418 -35
rect 420 -37 441 -35
rect 443 -37 444 -35
rect 539 -35 540 -33
rect 542 -35 544 -33
rect 539 -36 544 -35
rect 569 -33 622 -32
rect 569 -35 570 -33
rect 572 -35 622 -33
rect 569 -36 622 -35
rect 711 -35 764 -32
rect 711 -36 793 -35
rect 417 -38 444 -37
rect 618 -38 622 -36
rect 760 -38 790 -36
rect 792 -38 793 -36
rect 618 -39 671 -38
rect 760 -39 793 -38
rect 488 -41 614 -40
rect 488 -43 489 -41
rect 491 -43 611 -41
rect 613 -43 614 -41
rect 618 -41 668 -39
rect 670 -41 671 -39
rect 618 -42 671 -41
rect 718 -41 722 -40
rect 488 -44 614 -43
rect 718 -43 719 -41
rect 721 -43 722 -41
rect 718 -48 722 -43
rect 766 -44 770 -43
rect 766 -46 767 -44
rect 769 -46 770 -44
rect 660 -49 723 -48
rect 660 -51 661 -49
rect 663 -51 723 -49
rect 660 -52 723 -51
rect 766 -50 770 -46
rect 766 -52 767 -50
rect 769 -52 770 -50
rect 766 -53 770 -52
rect 761 -65 769 -62
rect 761 -67 762 -65
rect 764 -67 766 -65
rect 768 -67 769 -65
rect 761 -70 769 -67
rect 660 -81 721 -80
rect 660 -83 661 -81
rect 663 -83 721 -81
rect 660 -84 721 -83
rect 417 -89 439 -88
rect 417 -91 418 -89
rect 420 -91 436 -89
rect 438 -91 439 -89
rect 417 -92 439 -91
rect 488 -89 614 -88
rect 488 -91 489 -89
rect 491 -91 611 -89
rect 613 -91 614 -89
rect 488 -92 614 -91
rect 717 -89 721 -84
rect 717 -91 718 -89
rect 720 -91 721 -89
rect 717 -92 721 -91
rect 766 -89 770 -88
rect 766 -91 767 -89
rect 769 -91 770 -89
rect 699 -93 707 -92
rect 699 -95 700 -93
rect 702 -95 704 -93
rect 706 -95 707 -93
rect 699 -96 707 -95
rect 766 -93 770 -91
rect 766 -95 767 -93
rect 769 -95 770 -93
rect 766 -96 770 -95
rect 489 -97 542 -96
rect 489 -99 490 -97
rect 492 -99 539 -97
rect 541 -99 542 -97
rect 489 -100 542 -99
rect 569 -97 672 -96
rect 569 -99 570 -97
rect 572 -99 668 -97
rect 670 -99 672 -97
rect 569 -100 672 -99
rect 480 -105 529 -104
rect 480 -107 481 -105
rect 483 -107 526 -105
rect 528 -107 529 -105
rect 480 -108 529 -107
rect 627 -105 695 -104
rect 627 -107 628 -105
rect 630 -107 692 -105
rect 694 -107 695 -105
rect 627 -108 695 -107
rect 743 -105 753 -103
rect 743 -107 745 -105
rect 747 -107 750 -105
rect 752 -107 753 -105
rect 743 -108 753 -107
rect 800 -105 809 -104
rect 800 -107 801 -105
rect 803 -107 806 -105
rect 808 -107 809 -105
rect 800 -108 809 -107
rect 830 -108 834 -107
rect 579 -110 623 -109
rect 579 -112 580 -110
rect 582 -112 623 -110
rect 830 -110 831 -108
rect 833 -110 834 -108
rect 830 -112 834 -110
rect 579 -113 623 -112
rect 716 -113 779 -112
rect 619 -114 671 -113
rect 619 -116 668 -114
rect 670 -116 671 -114
rect 716 -115 719 -113
rect 721 -115 730 -113
rect 732 -115 775 -113
rect 777 -115 779 -113
rect 830 -114 831 -112
rect 833 -114 834 -112
rect 830 -115 834 -114
rect 716 -116 779 -115
rect 619 -117 671 -116
rect 309 -119 429 -118
rect 309 -121 310 -119
rect 312 -121 425 -119
rect 427 -121 429 -119
rect 309 -122 429 -121
rect 528 -126 748 -125
rect 528 -128 529 -126
rect 531 -128 744 -126
rect 746 -128 748 -126
rect 528 -129 748 -128
rect 834 -137 838 -136
rect 834 -139 835 -137
rect 837 -139 838 -137
rect 834 -140 838 -139
rect 834 -142 835 -140
rect 837 -142 838 -140
rect 834 -143 838 -142
rect 261 -148 751 -147
rect 261 -150 262 -148
rect 264 -150 748 -148
rect 750 -150 751 -148
rect 261 -151 751 -150
rect 50 -159 429 -158
rect 50 -161 51 -159
rect 53 -161 426 -159
rect 428 -161 429 -159
rect 50 -163 429 -161
rect 717 -161 779 -160
rect 717 -163 718 -161
rect 720 -163 730 -161
rect 732 -163 776 -161
rect 778 -163 779 -161
rect 579 -164 671 -163
rect 717 -164 779 -163
rect 579 -166 580 -164
rect 582 -166 668 -164
rect 670 -166 671 -164
rect 579 -167 671 -166
rect 830 -165 834 -164
rect 830 -167 831 -165
rect 833 -167 834 -165
rect 830 -168 834 -167
rect 480 -169 524 -168
rect 480 -171 481 -169
rect 483 -171 521 -169
rect 523 -171 524 -169
rect 744 -169 751 -168
rect 744 -171 745 -169
rect 747 -171 748 -169
rect 750 -171 751 -169
rect 480 -172 524 -171
rect 627 -172 707 -171
rect 744 -172 751 -171
rect 766 -169 770 -168
rect 766 -171 767 -169
rect 769 -171 770 -169
rect 766 -172 770 -171
rect 627 -174 628 -172
rect 630 -174 704 -172
rect 706 -174 707 -172
rect 627 -175 707 -174
rect 766 -174 767 -172
rect 769 -174 770 -172
rect 806 -170 814 -169
rect 806 -172 807 -170
rect 809 -172 811 -170
rect 813 -172 814 -170
rect 830 -170 831 -168
rect 833 -170 834 -168
rect 830 -171 834 -170
rect 806 -173 814 -172
rect 766 -176 770 -174
rect 507 -177 543 -176
rect 507 -179 508 -177
rect 510 -179 540 -177
rect 542 -179 543 -177
rect 507 -180 543 -179
rect 569 -177 622 -176
rect 569 -179 570 -177
rect 572 -179 622 -177
rect 569 -180 622 -179
rect 618 -182 622 -180
rect 691 -182 703 -181
rect 618 -183 671 -182
rect 488 -185 614 -184
rect 417 -186 437 -185
rect 417 -188 418 -186
rect 420 -188 434 -186
rect 436 -188 437 -186
rect 488 -187 489 -185
rect 491 -187 611 -185
rect 613 -187 614 -185
rect 618 -185 668 -183
rect 670 -185 671 -183
rect 691 -184 692 -182
rect 694 -184 700 -182
rect 702 -184 703 -182
rect 691 -185 703 -184
rect 717 -185 721 -184
rect 618 -186 671 -185
rect 488 -188 614 -187
rect 717 -187 718 -185
rect 720 -187 721 -185
rect 417 -189 437 -188
rect 717 -192 721 -187
rect 660 -193 721 -192
rect 660 -195 661 -193
rect 663 -195 721 -193
rect 660 -196 721 -195
rect 764 -209 772 -206
rect 764 -211 765 -209
rect 767 -211 769 -209
rect 771 -211 772 -209
rect 764 -214 772 -211
rect 660 -225 721 -224
rect 660 -227 661 -225
rect 663 -227 721 -225
rect 660 -228 721 -227
rect 417 -232 438 -231
rect 417 -234 418 -232
rect 420 -234 435 -232
rect 437 -234 438 -232
rect 417 -235 438 -234
rect 488 -233 614 -232
rect 488 -235 489 -233
rect 491 -235 611 -233
rect 613 -235 614 -233
rect 488 -236 614 -235
rect 717 -233 721 -228
rect 717 -235 718 -233
rect 720 -235 721 -233
rect 717 -236 721 -235
rect 699 -237 707 -236
rect 699 -239 700 -237
rect 702 -239 704 -237
rect 706 -239 707 -237
rect 699 -240 707 -239
rect 463 -241 543 -240
rect 463 -243 464 -241
rect 466 -243 540 -241
rect 542 -243 543 -241
rect 463 -244 543 -243
rect 569 -241 672 -240
rect 569 -243 570 -241
rect 572 -243 668 -241
rect 670 -243 672 -241
rect 569 -244 672 -243
rect 480 -249 534 -248
rect 480 -251 481 -249
rect 483 -251 531 -249
rect 533 -251 534 -249
rect 480 -252 534 -251
rect 617 -249 625 -248
rect 617 -251 618 -249
rect 620 -251 622 -249
rect 624 -251 625 -249
rect 617 -252 625 -251
rect 745 -249 752 -248
rect 745 -251 746 -249
rect 748 -251 749 -249
rect 751 -251 752 -249
rect 745 -252 752 -251
rect 766 -249 770 -248
rect 766 -251 767 -249
rect 769 -251 770 -249
rect 766 -253 770 -251
rect 813 -249 824 -248
rect 813 -251 814 -249
rect 816 -251 821 -249
rect 823 -251 824 -249
rect 813 -252 824 -251
rect 830 -249 834 -248
rect 830 -251 831 -249
rect 833 -251 834 -249
rect 579 -254 613 -253
rect 0 -255 429 -254
rect 0 -257 1 -255
rect 3 -257 426 -255
rect 428 -257 429 -255
rect 579 -256 580 -254
rect 582 -256 613 -254
rect 579 -257 613 -256
rect 632 -254 671 -253
rect 632 -256 668 -254
rect 670 -256 671 -254
rect 766 -255 767 -253
rect 769 -255 770 -253
rect 766 -256 770 -255
rect 830 -253 834 -251
rect 830 -255 831 -253
rect 833 -255 834 -253
rect 830 -256 834 -255
rect 632 -257 671 -256
rect 0 -258 429 -257
rect 608 -261 636 -257
rect 710 -266 779 -265
rect 710 -268 712 -266
rect 714 -268 730 -266
rect 732 -268 776 -266
rect 778 -268 779 -266
rect 417 -269 621 -268
rect 710 -269 779 -268
rect 417 -271 418 -269
rect 420 -271 618 -269
rect 620 -271 621 -269
rect 417 -272 621 -271
rect 528 -279 537 -278
rect 460 -280 469 -279
rect 460 -282 461 -280
rect 463 -282 466 -280
rect 468 -282 469 -280
rect 460 -283 469 -282
rect 528 -281 529 -279
rect 531 -280 537 -279
rect 531 -281 534 -280
rect 528 -282 534 -281
rect 536 -282 537 -280
rect 528 -283 537 -282
rect 611 -279 620 -278
rect 611 -281 612 -279
rect 614 -280 620 -279
rect 614 -281 617 -280
rect 611 -282 617 -281
rect 619 -282 620 -280
rect 611 -283 620 -282
rect 708 -279 717 -278
rect 708 -281 709 -279
rect 711 -280 717 -279
rect 711 -281 714 -280
rect 708 -282 714 -281
rect 716 -282 717 -280
rect 708 -283 717 -282
rect 772 -279 781 -278
rect 772 -281 773 -279
rect 775 -280 781 -279
rect 775 -281 778 -280
rect 772 -282 778 -281
rect 780 -282 781 -280
rect 772 -283 781 -282
<< alu3 >>
rect 30 305 34 306
rect 30 303 31 305
rect 33 303 34 305
rect 30 294 34 303
rect 30 292 31 294
rect 33 292 34 294
rect 30 291 34 292
rect 163 305 167 306
rect 163 303 164 305
rect 166 303 167 305
rect 163 294 167 303
rect 163 292 164 294
rect 166 292 167 294
rect 163 291 167 292
rect 403 305 407 306
rect 403 303 404 305
rect 406 303 407 305
rect 403 294 407 303
rect 403 292 404 294
rect 406 292 407 294
rect 403 291 407 292
rect 588 305 592 306
rect 588 303 589 305
rect 591 303 592 305
rect 588 294 592 303
rect 588 292 589 294
rect 591 292 592 294
rect 588 291 592 292
rect 780 305 784 306
rect 780 303 781 305
rect 783 303 784 305
rect 780 294 784 303
rect 780 292 781 294
rect 783 292 784 294
rect 780 291 784 292
rect 30 285 34 286
rect 30 283 31 285
rect 33 283 34 285
rect 0 266 4 267
rect 0 264 1 266
rect 3 264 4 266
rect 0 195 4 264
rect 20 246 24 247
rect 20 244 21 246
rect 23 244 24 246
rect 20 223 24 244
rect 20 221 21 223
rect 23 221 24 223
rect 20 220 24 221
rect 0 193 1 195
rect 3 193 4 195
rect -10 138 -6 139
rect -10 136 -9 138
rect -7 136 -6 138
rect -10 135 -6 136
rect -10 133 -9 135
rect -7 133 -6 135
rect -10 132 -6 133
rect 0 122 4 193
rect 14 174 18 176
rect 14 172 15 174
rect 17 172 18 174
rect 14 151 18 172
rect 14 149 15 151
rect 17 149 18 151
rect 14 148 18 149
rect 0 120 1 122
rect 3 120 4 122
rect 0 35 4 120
rect 22 103 26 104
rect 22 101 23 103
rect 25 101 26 103
rect 22 79 26 101
rect 22 77 23 79
rect 25 77 26 79
rect 22 76 26 77
rect 30 55 34 283
rect 52 285 56 286
rect 52 283 53 285
rect 55 283 56 285
rect 52 272 56 283
rect 52 270 53 272
rect 55 270 56 272
rect 52 269 56 270
rect 304 285 308 286
rect 304 283 305 285
rect 307 283 308 285
rect 304 272 308 283
rect 304 270 305 272
rect 307 270 308 272
rect 304 269 308 270
rect 463 285 467 286
rect 463 283 464 285
rect 466 283 467 285
rect 210 263 214 264
rect 210 261 211 263
rect 213 261 214 263
rect 30 53 31 55
rect 33 53 34 55
rect 30 52 34 53
rect 42 249 46 250
rect 42 247 43 249
rect 45 247 46 249
rect 42 175 46 247
rect 210 226 214 261
rect 332 263 336 264
rect 332 261 333 263
rect 335 261 336 263
rect 301 251 305 252
rect 301 249 302 251
rect 304 249 305 251
rect 210 224 211 226
rect 213 224 214 226
rect 61 223 65 224
rect 210 223 214 224
rect 261 244 265 245
rect 261 242 262 244
rect 264 242 265 244
rect 61 221 62 223
rect 64 221 65 223
rect 61 197 65 221
rect 61 195 62 197
rect 64 195 65 197
rect 61 194 65 195
rect 42 173 43 175
rect 45 173 46 175
rect 42 106 46 173
rect 63 151 67 152
rect 63 149 64 151
rect 66 149 67 151
rect 63 128 67 149
rect 63 126 64 128
rect 66 126 67 128
rect 63 125 67 126
rect 42 104 43 106
rect 45 104 46 106
rect 42 51 46 104
rect 61 79 65 80
rect 61 77 62 79
rect 64 77 65 79
rect 61 56 65 77
rect 61 54 62 56
rect 64 54 65 56
rect 61 53 65 54
rect 126 76 130 77
rect 126 74 127 76
rect 129 74 130 76
rect 42 50 54 51
rect 42 48 43 50
rect 45 48 54 50
rect 42 47 54 48
rect 0 33 1 35
rect 3 33 4 35
rect 0 -49 4 33
rect 38 22 42 23
rect 38 20 39 22
rect 41 20 42 22
rect 19 11 24 12
rect 19 9 20 11
rect 22 9 24 11
rect 19 8 24 9
rect 19 6 20 8
rect 22 6 24 8
rect 19 5 24 6
rect 38 4 42 20
rect 38 2 39 4
rect 41 2 42 4
rect 38 1 42 2
rect 0 -51 1 -49
rect 3 -51 4 -49
rect 0 -255 4 -51
rect 50 -39 54 47
rect 126 39 130 74
rect 126 37 127 39
rect 129 37 130 39
rect 126 36 130 37
rect 50 -41 51 -39
rect 53 -41 54 -39
rect 50 -159 54 -41
rect 261 -148 265 242
rect 289 223 293 224
rect 289 221 290 223
rect 292 221 293 223
rect 289 198 293 221
rect 289 196 290 198
rect 292 196 293 198
rect 289 195 293 196
rect 301 186 305 249
rect 301 184 302 186
rect 304 184 305 186
rect 301 183 305 184
rect 309 249 313 250
rect 309 247 310 249
rect 312 247 313 249
rect 309 175 313 247
rect 332 207 336 261
rect 332 205 333 207
rect 335 205 336 207
rect 332 204 336 205
rect 309 173 310 175
rect 312 173 313 175
rect 298 151 302 152
rect 298 149 299 151
rect 301 149 302 151
rect 298 124 302 149
rect 298 122 299 124
rect 301 122 302 124
rect 298 121 302 122
rect 301 107 305 108
rect 301 105 302 107
rect 304 105 305 107
rect 289 79 293 80
rect 289 77 290 79
rect 292 77 293 79
rect 289 52 293 77
rect 289 50 290 52
rect 292 50 293 52
rect 289 49 293 50
rect 301 42 305 105
rect 301 40 302 42
rect 304 40 305 42
rect 301 39 305 40
rect 309 106 313 173
rect 309 104 310 106
rect 312 104 313 106
rect 309 34 313 104
rect 320 183 324 184
rect 320 181 321 183
rect 323 181 324 183
rect 320 95 324 181
rect 320 93 321 95
rect 323 93 324 95
rect 320 92 324 93
rect 333 119 337 120
rect 333 117 334 119
rect 336 117 337 119
rect 333 63 337 117
rect 333 61 334 63
rect 336 61 337 63
rect 333 60 337 61
rect 309 32 310 34
rect 312 32 313 34
rect 309 -26 313 32
rect 393 39 397 40
rect 393 37 394 39
rect 396 37 397 39
rect 393 23 397 37
rect 393 21 394 23
rect 396 21 397 23
rect 393 19 397 21
rect 404 4 408 5
rect 404 2 405 4
rect 407 2 408 4
rect 389 -8 393 -7
rect 389 -10 390 -8
rect 392 -10 393 -8
rect 389 -12 393 -10
rect 389 -14 390 -12
rect 392 -14 393 -12
rect 389 -15 393 -14
rect 309 -28 310 -26
rect 312 -28 313 -26
rect 309 -119 313 -28
rect 309 -121 310 -119
rect 312 -121 313 -119
rect 309 -122 313 -121
rect 261 -150 262 -148
rect 264 -150 265 -148
rect 261 -151 265 -150
rect 50 -161 51 -159
rect 53 -161 54 -159
rect 50 -163 54 -161
rect 0 -257 1 -255
rect 3 -257 4 -255
rect 0 -258 4 -257
rect 404 -258 408 2
rect 404 -260 405 -258
rect 407 -260 408 -258
rect 404 -261 408 -260
rect 417 -35 421 -34
rect 417 -37 418 -35
rect 420 -37 421 -35
rect 417 -89 421 -37
rect 417 -91 418 -89
rect 420 -91 421 -89
rect 417 -186 421 -91
rect 417 -188 418 -186
rect 420 -188 421 -186
rect 417 -232 421 -188
rect 417 -234 418 -232
rect 420 -234 421 -232
rect 417 -269 421 -234
rect 463 -241 467 283
rect 573 285 577 286
rect 573 283 574 285
rect 576 283 577 285
rect 573 272 577 283
rect 573 270 574 272
rect 576 270 577 272
rect 573 269 577 270
rect 477 263 481 264
rect 477 261 478 263
rect 480 261 481 263
rect 477 226 481 261
rect 599 263 603 264
rect 599 261 600 263
rect 602 261 603 263
rect 568 251 572 252
rect 568 249 569 251
rect 571 249 572 251
rect 477 224 478 226
rect 480 224 481 226
rect 528 245 532 246
rect 528 243 529 245
rect 531 243 532 245
rect 477 223 481 224
rect 507 223 511 224
rect 507 221 508 223
rect 510 221 511 223
rect 489 151 493 152
rect 489 149 490 151
rect 492 149 493 151
rect 489 -97 493 149
rect 489 -99 490 -97
rect 492 -99 493 -97
rect 489 -100 493 -99
rect 507 -177 511 221
rect 528 -126 532 243
rect 554 223 558 224
rect 554 221 555 223
rect 557 221 558 223
rect 554 196 558 221
rect 554 194 555 196
rect 557 194 558 196
rect 554 193 558 194
rect 568 186 572 249
rect 568 184 569 186
rect 571 184 572 186
rect 568 183 572 184
rect 576 249 580 250
rect 576 247 577 249
rect 579 247 580 249
rect 576 175 580 247
rect 599 207 603 261
rect 744 263 748 264
rect 744 261 745 263
rect 747 261 748 263
rect 744 226 748 261
rect 835 251 839 252
rect 835 249 836 251
rect 838 249 839 251
rect 744 224 745 226
rect 747 224 748 226
rect 744 223 748 224
rect 754 245 758 246
rect 754 243 755 245
rect 757 243 758 245
rect 599 205 600 207
rect 602 205 603 207
rect 599 204 603 205
rect 576 173 577 175
rect 579 173 580 175
rect 567 151 571 152
rect 567 149 568 151
rect 570 149 571 151
rect 567 128 571 149
rect 567 126 568 128
rect 570 126 571 128
rect 567 125 571 126
rect 568 107 572 108
rect 568 105 569 107
rect 571 105 572 107
rect 540 79 544 80
rect 540 77 541 79
rect 543 77 544 79
rect 540 -27 544 77
rect 551 79 555 80
rect 551 77 552 79
rect 554 77 555 79
rect 551 53 555 77
rect 551 51 552 53
rect 554 51 555 53
rect 551 50 555 51
rect 568 42 572 105
rect 568 40 569 42
rect 571 40 572 42
rect 568 39 572 40
rect 576 106 580 173
rect 576 104 577 106
rect 579 104 580 106
rect 576 34 580 104
rect 588 183 592 184
rect 588 181 589 183
rect 591 181 592 183
rect 588 95 592 181
rect 588 93 589 95
rect 591 93 592 95
rect 588 92 592 93
rect 599 119 604 120
rect 599 117 600 119
rect 602 117 604 119
rect 599 64 604 117
rect 599 62 601 64
rect 603 62 604 64
rect 599 60 604 62
rect 576 32 577 34
rect 579 32 580 34
rect 576 -8 580 32
rect 660 39 664 40
rect 660 37 661 39
rect 663 37 664 39
rect 660 22 664 37
rect 660 20 661 22
rect 663 20 664 22
rect 660 19 664 20
rect 576 -10 577 -8
rect 579 -10 580 -8
rect 576 -11 580 -10
rect 729 -17 733 -16
rect 729 -19 730 -17
rect 732 -19 733 -17
rect 540 -29 541 -27
rect 543 -29 544 -27
rect 540 -30 544 -29
rect 703 -28 707 -27
rect 703 -30 704 -28
rect 706 -30 707 -28
rect 703 -93 707 -30
rect 703 -95 704 -93
rect 706 -95 707 -93
rect 703 -96 707 -95
rect 528 -128 529 -126
rect 531 -128 532 -126
rect 528 -129 532 -128
rect 691 -105 695 -104
rect 691 -107 692 -105
rect 694 -107 695 -105
rect 507 -179 508 -177
rect 510 -179 511 -177
rect 507 -180 511 -179
rect 691 -182 695 -107
rect 729 -113 733 -19
rect 754 -23 758 243
rect 772 223 780 226
rect 772 221 773 223
rect 775 221 777 223
rect 779 221 780 223
rect 772 218 780 221
rect 788 208 792 209
rect 788 206 789 208
rect 791 206 792 208
rect 766 79 774 82
rect 766 77 767 79
rect 769 77 771 79
rect 773 77 774 79
rect 766 74 774 77
rect 750 -25 758 -23
rect 750 -27 751 -25
rect 753 -27 758 -25
rect 750 -28 758 -27
rect 788 -26 792 206
rect 835 186 839 249
rect 835 184 836 186
rect 838 184 839 186
rect 835 183 839 184
rect 833 154 848 155
rect 833 152 834 154
rect 836 152 845 154
rect 847 152 848 154
rect 833 151 848 152
rect 835 107 839 108
rect 835 105 836 107
rect 838 105 839 107
rect 788 -28 789 -26
rect 791 -28 792 -26
rect 788 -29 792 -28
rect 800 95 804 96
rect 800 93 801 95
rect 803 93 804 95
rect 766 -40 770 -39
rect 766 -42 767 -40
rect 769 -42 770 -40
rect 766 -44 770 -42
rect 766 -46 767 -44
rect 769 -46 770 -44
rect 766 -47 770 -46
rect 765 -65 773 -62
rect 765 -67 766 -65
rect 768 -67 770 -65
rect 772 -67 773 -65
rect 765 -70 773 -67
rect 766 -93 770 -92
rect 766 -95 767 -93
rect 769 -95 770 -93
rect 766 -97 770 -95
rect 766 -99 767 -97
rect 769 -99 770 -97
rect 766 -100 770 -99
rect 729 -115 730 -113
rect 732 -115 733 -113
rect 729 -161 733 -115
rect 743 -105 748 -103
rect 743 -107 745 -105
rect 747 -107 748 -105
rect 743 -126 748 -107
rect 800 -105 804 93
rect 800 -107 801 -105
rect 803 -107 804 -105
rect 800 -108 804 -107
rect 810 63 814 64
rect 810 61 811 63
rect 813 61 814 63
rect 743 -128 744 -126
rect 746 -128 748 -126
rect 743 -129 748 -128
rect 729 -163 730 -161
rect 732 -163 733 -161
rect 691 -184 692 -182
rect 694 -184 695 -182
rect 691 -185 695 -184
rect 703 -172 707 -171
rect 703 -174 704 -172
rect 706 -174 707 -172
rect 703 -237 707 -174
rect 703 -239 704 -237
rect 706 -239 707 -237
rect 703 -240 707 -239
rect 463 -243 464 -241
rect 466 -243 467 -241
rect 463 -244 467 -243
rect 417 -271 418 -269
rect 420 -271 421 -269
rect 417 -272 421 -271
rect 617 -249 621 -248
rect 617 -251 618 -249
rect 620 -251 621 -249
rect 617 -269 621 -251
rect 617 -271 618 -269
rect 620 -271 621 -269
rect 617 -272 621 -271
rect 729 -266 733 -163
rect 747 -148 751 -147
rect 747 -150 748 -148
rect 750 -150 751 -148
rect 747 -169 751 -150
rect 747 -171 748 -169
rect 750 -171 751 -169
rect 810 -170 814 61
rect 835 42 839 105
rect 835 40 836 42
rect 838 40 839 42
rect 835 39 839 40
rect 747 -172 751 -171
rect 766 -172 770 -171
rect 766 -174 767 -172
rect 769 -174 770 -172
rect 810 -172 811 -170
rect 813 -172 814 -170
rect 810 -173 814 -172
rect 820 23 824 24
rect 820 21 821 23
rect 823 21 824 23
rect 766 -175 770 -174
rect 766 -177 767 -175
rect 769 -177 770 -175
rect 766 -178 770 -177
rect 767 -209 780 -206
rect 767 -211 769 -209
rect 771 -211 773 -209
rect 775 -211 780 -209
rect 767 -214 780 -211
rect 766 -245 770 -244
rect 766 -247 767 -245
rect 769 -247 770 -245
rect 745 -249 749 -248
rect 745 -251 746 -249
rect 748 -251 749 -249
rect 745 -258 749 -251
rect 766 -249 770 -247
rect 766 -251 767 -249
rect 769 -251 770 -249
rect 766 -252 770 -251
rect 820 -249 824 21
rect 832 10 847 11
rect 832 8 833 10
rect 835 8 844 10
rect 846 8 847 10
rect 832 7 847 8
rect 861 1 865 2
rect 861 -1 862 1
rect 864 -1 865 1
rect 830 -20 834 -19
rect 830 -22 831 -20
rect 833 -22 834 -20
rect 830 -23 834 -22
rect 830 -25 831 -23
rect 833 -25 834 -23
rect 830 -26 834 -25
rect 830 -112 834 -111
rect 830 -114 831 -112
rect 833 -114 834 -112
rect 830 -116 834 -114
rect 830 -118 831 -116
rect 833 -118 834 -116
rect 830 -119 834 -118
rect 834 -137 849 -136
rect 834 -139 835 -137
rect 837 -139 846 -137
rect 848 -139 849 -137
rect 834 -140 849 -139
rect 830 -162 834 -161
rect 830 -164 831 -162
rect 833 -164 834 -162
rect 830 -165 834 -164
rect 830 -167 831 -165
rect 833 -167 834 -165
rect 830 -168 834 -167
rect 820 -251 821 -249
rect 823 -251 824 -249
rect 820 -252 824 -251
rect 745 -260 746 -258
rect 748 -260 749 -258
rect 830 -253 834 -252
rect 830 -255 831 -253
rect 833 -255 834 -253
rect 830 -257 834 -255
rect 830 -259 831 -257
rect 833 -259 834 -257
rect 830 -260 834 -259
rect 861 -257 865 -1
rect 869 -7 873 -6
rect 869 -9 870 -7
rect 872 -9 873 -7
rect 869 -162 873 -9
rect 877 -15 881 -14
rect 877 -17 878 -15
rect 880 -17 881 -15
rect 877 -116 881 -17
rect 877 -118 878 -116
rect 880 -118 881 -116
rect 877 -119 881 -118
rect 869 -164 870 -162
rect 872 -164 873 -162
rect 869 -165 873 -164
rect 861 -259 862 -257
rect 864 -259 865 -257
rect 861 -260 865 -259
rect 745 -261 749 -260
rect 729 -268 730 -266
rect 732 -268 733 -266
rect 729 -271 733 -268
rect 729 -273 730 -271
rect 732 -273 733 -271
rect 729 -274 733 -273
rect 465 -280 469 -279
rect 465 -282 466 -280
rect 468 -282 469 -280
rect 465 -291 469 -282
rect 465 -293 466 -291
rect 468 -293 469 -291
rect 465 -294 469 -293
rect 533 -280 537 -279
rect 533 -282 534 -280
rect 536 -282 537 -280
rect 533 -291 537 -282
rect 533 -293 534 -291
rect 536 -293 537 -291
rect 533 -294 537 -293
rect 616 -280 620 -279
rect 616 -282 617 -280
rect 619 -282 620 -280
rect 616 -291 620 -282
rect 616 -293 617 -291
rect 619 -293 620 -291
rect 616 -294 620 -293
rect 713 -280 717 -279
rect 713 -282 714 -280
rect 716 -282 717 -280
rect 713 -291 717 -282
rect 713 -293 714 -291
rect 716 -293 717 -291
rect 713 -294 717 -293
rect 777 -280 781 -279
rect 777 -282 778 -280
rect 780 -282 781 -280
rect 777 -291 781 -282
rect 777 -293 778 -291
rect 780 -293 781 -291
rect 777 -294 781 -293
<< alu4 >>
rect 27 305 34 306
rect 27 303 28 305
rect 30 303 31 305
rect 33 303 34 305
rect 27 302 34 303
rect 160 305 167 306
rect 160 303 161 305
rect 163 303 164 305
rect 166 303 167 305
rect 160 302 167 303
rect 400 305 407 306
rect 400 303 401 305
rect 403 303 404 305
rect 406 303 407 305
rect 400 302 407 303
rect 585 305 592 306
rect 585 303 586 305
rect 588 303 589 305
rect 591 303 592 305
rect 585 302 592 303
rect 777 305 784 306
rect 777 303 778 305
rect 780 303 781 305
rect 783 303 784 305
rect 777 302 784 303
rect -39 286 2 287
rect -39 285 577 286
rect -39 283 31 285
rect 33 283 53 285
rect 55 283 305 285
rect 307 283 464 285
rect 466 283 574 285
rect 576 283 577 285
rect -39 282 577 283
rect -39 234 -34 282
rect -49 229 -34 234
rect -49 224 8 225
rect -49 223 558 224
rect -49 221 21 223
rect 23 221 62 223
rect 64 221 290 223
rect 292 221 508 223
rect 510 221 555 223
rect 557 221 558 223
rect -49 220 558 221
rect 776 223 785 226
rect 776 221 777 223
rect 779 221 782 223
rect 784 221 785 223
rect 776 218 785 221
rect -49 208 -25 213
rect -49 197 -36 202
rect -42 81 -36 197
rect -31 153 -25 208
rect 844 154 848 155
rect -31 152 10 153
rect 844 152 845 154
rect 847 152 848 154
rect -31 151 571 152
rect -31 149 15 151
rect 17 149 64 151
rect 66 149 299 151
rect 301 149 490 151
rect 492 149 568 151
rect 570 149 571 151
rect -31 148 571 149
rect 844 151 848 152
rect 844 149 845 151
rect 847 149 848 151
rect 844 148 848 149
rect -10 141 -6 142
rect -10 139 -9 141
rect -7 139 -6 141
rect -10 138 -6 139
rect -10 136 -9 138
rect -7 136 -6 138
rect -10 135 -6 136
rect -42 80 2 81
rect -42 79 556 80
rect -42 77 23 79
rect 25 77 62 79
rect 64 77 290 79
rect 292 77 541 79
rect 543 77 552 79
rect 554 77 556 79
rect -42 76 556 77
rect 770 79 778 82
rect 770 77 771 79
rect 773 77 775 79
rect 777 77 778 79
rect 770 74 778 77
rect -10 11 24 12
rect -10 9 -9 11
rect -7 9 20 11
rect 22 9 24 11
rect -10 8 24 9
rect 843 10 847 11
rect 843 8 844 10
rect 846 8 847 10
rect 843 7 847 8
rect 843 5 844 7
rect 846 5 847 7
rect 843 4 847 5
rect 861 1 908 2
rect 861 -1 862 1
rect 864 -1 908 1
rect 861 -2 908 -1
rect 869 -7 908 -6
rect 869 -9 870 -7
rect 872 -9 908 -7
rect 869 -10 908 -9
rect -73 -12 393 -11
rect -73 -14 390 -12
rect 392 -14 393 -12
rect -73 -16 393 -14
rect 877 -15 908 -14
rect 877 -17 878 -15
rect 880 -17 908 -15
rect 877 -18 908 -17
rect 830 -23 908 -22
rect 830 -25 831 -23
rect 833 -25 908 -23
rect -73 -26 313 -25
rect 830 -26 908 -25
rect -73 -28 310 -26
rect 312 -28 313 -26
rect -73 -29 313 -28
rect -73 -39 54 -38
rect -73 -41 51 -39
rect 53 -41 54 -39
rect -73 -42 54 -41
rect 766 -40 908 -39
rect 766 -42 767 -40
rect 769 -42 908 -40
rect 766 -43 908 -42
rect -73 -49 4 -48
rect -73 -51 1 -49
rect 3 -51 4 -49
rect -73 -52 4 -51
rect 882 -51 908 -47
rect 769 -65 777 -62
rect 769 -67 770 -65
rect 772 -67 774 -65
rect 776 -67 777 -65
rect 769 -70 777 -67
rect 882 -96 886 -51
rect 766 -97 886 -96
rect 766 -99 767 -97
rect 769 -99 886 -97
rect 766 -100 886 -99
rect 890 -59 908 -55
rect 830 -116 881 -115
rect 830 -118 831 -116
rect 833 -118 878 -116
rect 880 -118 881 -116
rect 830 -119 881 -118
rect 845 -137 849 -136
rect 845 -139 846 -137
rect 848 -139 849 -137
rect 845 -141 849 -139
rect 845 -143 846 -141
rect 848 -143 849 -141
rect 845 -144 849 -143
rect 830 -162 873 -161
rect 830 -164 831 -162
rect 833 -164 870 -162
rect 872 -164 873 -162
rect 830 -165 873 -164
rect 890 -174 894 -59
rect 766 -175 894 -174
rect 766 -177 767 -175
rect 769 -177 894 -175
rect 766 -178 894 -177
rect 901 -67 908 -63
rect 772 -209 781 -208
rect 772 -211 773 -209
rect 775 -211 778 -209
rect 780 -211 781 -209
rect 772 -212 781 -211
rect 901 -244 905 -67
rect 766 -245 905 -244
rect 766 -247 767 -245
rect 769 -247 905 -245
rect 766 -248 905 -247
rect 830 -257 865 -256
rect 404 -258 749 -257
rect 404 -260 405 -258
rect 407 -260 746 -258
rect 748 -260 749 -258
rect 830 -259 831 -257
rect 833 -259 862 -257
rect 864 -259 865 -257
rect 830 -260 865 -259
rect 404 -261 749 -260
rect -49 -271 733 -270
rect -49 -273 730 -271
rect 732 -273 733 -271
rect -49 -275 733 -273
rect 462 -291 469 -290
rect 462 -293 463 -291
rect 465 -293 466 -291
rect 468 -293 469 -291
rect 462 -294 469 -293
rect 530 -291 537 -290
rect 530 -293 531 -291
rect 533 -293 534 -291
rect 536 -293 537 -291
rect 530 -294 537 -293
rect 613 -291 620 -290
rect 613 -293 614 -291
rect 616 -293 617 -291
rect 619 -293 620 -291
rect 613 -294 620 -293
rect 710 -291 717 -290
rect 710 -293 711 -291
rect 713 -293 714 -291
rect 716 -293 717 -291
rect 710 -294 717 -293
rect 774 -291 781 -290
rect 774 -293 775 -291
rect 777 -293 778 -291
rect 780 -293 781 -291
rect 774 -294 781 -293
<< alu5 >>
rect -12 305 851 308
rect -12 303 28 305
rect 30 303 161 305
rect 163 303 401 305
rect 403 303 586 305
rect 588 303 778 305
rect 780 303 851 305
rect -12 300 851 303
rect -12 141 -4 300
rect 780 224 816 226
rect 780 223 810 224
rect 780 221 782 223
rect 784 221 810 223
rect 780 220 810 221
rect 814 220 816 224
rect 780 218 816 220
rect 843 155 851 300
rect 842 151 851 155
rect 842 149 845 151
rect 847 149 851 151
rect 842 146 851 149
rect -12 139 -9 141
rect -7 139 -4 141
rect -12 11 -4 139
rect 773 80 816 82
rect 773 79 810 80
rect 773 77 775 79
rect 777 77 810 79
rect 773 76 810 77
rect 814 76 816 80
rect 773 74 816 76
rect 843 11 851 146
rect -12 9 -9 11
rect -7 9 -4 11
rect -12 -292 -4 9
rect 841 7 851 11
rect 841 5 844 7
rect 846 5 851 7
rect 841 2 851 5
rect 772 -64 815 -62
rect 772 -65 809 -64
rect 772 -67 774 -65
rect 776 -67 809 -65
rect 772 -68 809 -67
rect 813 -68 815 -64
rect 772 -70 815 -68
rect 843 -141 851 2
rect 843 -143 846 -141
rect 848 -143 851 -141
rect 772 -208 815 -206
rect 772 -209 809 -208
rect 772 -211 778 -209
rect 780 -211 809 -209
rect 772 -212 809 -211
rect 813 -212 815 -208
rect 772 -214 815 -212
rect 460 -291 469 -288
rect 460 -292 463 -291
rect -12 -293 463 -292
rect 465 -292 469 -291
rect 528 -291 537 -288
rect 528 -292 531 -291
rect 465 -293 531 -292
rect 533 -292 537 -291
rect 611 -291 620 -288
rect 611 -292 614 -291
rect 533 -293 614 -292
rect 616 -292 620 -291
rect 708 -291 717 -288
rect 708 -292 711 -291
rect 616 -293 711 -292
rect 713 -292 717 -291
rect 772 -291 781 -288
rect 772 -292 775 -291
rect 713 -293 775 -292
rect 777 -292 781 -291
rect 843 -292 851 -143
rect 777 -293 851 -292
rect -12 -300 851 -293
<< alu6 >>
rect -25 309 860 318
rect -25 -302 -17 309
rect 806 226 819 228
rect 852 226 860 309
rect 806 224 860 226
rect 806 220 810 224
rect 814 220 860 224
rect 806 218 860 220
rect 806 216 819 218
rect 806 82 819 84
rect 852 82 860 218
rect 806 80 860 82
rect 806 76 810 80
rect 814 76 860 80
rect 806 74 860 76
rect 806 72 819 74
rect 805 -61 818 -60
rect 852 -61 860 74
rect 805 -64 860 -61
rect 805 -68 809 -64
rect 813 -68 860 -64
rect 805 -69 860 -68
rect 805 -72 818 -69
rect 805 -206 818 -204
rect 852 -206 860 -69
rect 805 -208 860 -206
rect 805 -212 809 -208
rect 813 -212 860 -208
rect 805 -214 860 -212
rect 805 -216 818 -214
rect 852 -302 860 -214
rect -25 -310 860 -302
<< ptie >>
rect 35 229 41 231
rect 35 227 37 229
rect 39 227 41 229
rect 35 225 41 227
rect 75 229 81 231
rect 75 227 77 229
rect 79 227 81 229
rect 75 225 81 227
rect 294 229 300 231
rect 294 227 296 229
rect 298 227 300 229
rect 294 225 300 227
rect 342 229 348 231
rect 342 227 344 229
rect 346 227 348 229
rect 342 225 348 227
rect 561 229 567 231
rect 561 227 563 229
rect 565 227 567 229
rect 561 225 567 227
rect 609 229 615 231
rect 609 227 611 229
rect 613 227 615 229
rect 609 225 615 227
rect 828 229 834 231
rect 828 227 830 229
rect 832 227 834 229
rect 828 225 834 227
rect 35 217 41 219
rect 35 215 37 217
rect 39 215 41 217
rect 35 213 41 215
rect 75 217 81 219
rect 75 215 77 217
rect 79 215 81 217
rect 75 213 81 215
rect 294 217 300 219
rect 294 215 296 217
rect 298 215 300 217
rect 294 213 300 215
rect 342 217 348 219
rect 342 215 344 217
rect 346 215 348 217
rect 342 213 348 215
rect 561 217 567 219
rect 561 215 563 217
rect 565 215 567 217
rect 561 213 567 215
rect 609 217 615 219
rect 609 215 611 217
rect 613 215 615 217
rect 609 213 615 215
rect 828 217 834 219
rect 828 215 830 217
rect 832 215 834 217
rect 828 213 834 215
rect 35 85 41 87
rect 35 83 37 85
rect 39 83 41 85
rect 35 81 41 83
rect 75 85 81 87
rect 75 83 77 85
rect 79 83 81 85
rect 75 81 81 83
rect 294 85 300 87
rect 294 83 296 85
rect 298 83 300 85
rect 294 81 300 83
rect 342 85 348 87
rect 342 83 344 85
rect 346 83 348 85
rect 342 81 348 83
rect 561 85 567 87
rect 561 83 563 85
rect 565 83 567 85
rect 561 81 567 83
rect 609 85 615 87
rect 609 83 611 85
rect 613 83 615 85
rect 609 81 615 83
rect 828 85 834 87
rect 828 83 830 85
rect 832 83 834 85
rect 828 81 834 83
rect 35 73 41 75
rect 35 71 37 73
rect 39 71 41 73
rect 35 69 41 71
rect 75 73 81 75
rect 75 71 77 73
rect 79 71 81 73
rect 75 69 81 71
rect 294 73 300 75
rect 294 71 296 73
rect 298 71 300 73
rect 294 69 300 71
rect 342 73 348 75
rect 342 71 344 73
rect 346 71 348 73
rect 342 69 348 71
rect 561 73 567 75
rect 561 71 563 73
rect 565 71 567 73
rect 561 69 567 71
rect 609 73 615 75
rect 609 71 611 73
rect 613 71 615 73
rect 609 69 615 71
rect 828 73 834 75
rect 828 71 830 73
rect 832 71 834 73
rect 828 69 834 71
rect 425 -59 431 -57
rect 425 -61 427 -59
rect 429 -61 431 -59
rect 425 -63 431 -61
rect 696 -59 702 -57
rect 696 -61 698 -59
rect 700 -61 702 -59
rect 696 -63 702 -61
rect 425 -71 431 -69
rect 425 -73 427 -71
rect 429 -73 431 -71
rect 425 -75 431 -73
rect 696 -71 702 -69
rect 696 -73 698 -71
rect 700 -73 702 -71
rect 696 -75 702 -73
rect 425 -203 431 -201
rect 425 -205 427 -203
rect 429 -205 431 -203
rect 425 -207 431 -205
rect 696 -203 702 -201
rect 696 -205 698 -203
rect 700 -205 702 -203
rect 696 -207 702 -205
rect 425 -215 431 -213
rect 425 -217 427 -215
rect 429 -217 431 -215
rect 425 -219 431 -217
rect 696 -215 702 -213
rect 696 -217 698 -215
rect 700 -217 702 -215
rect 696 -219 702 -217
<< ntie >>
rect 35 289 41 291
rect 35 287 37 289
rect 39 287 41 289
rect 35 285 41 287
rect 75 289 81 291
rect 75 287 77 289
rect 79 287 81 289
rect 75 285 81 287
rect 294 289 300 291
rect 294 287 296 289
rect 298 287 300 289
rect 294 285 300 287
rect 342 289 348 291
rect 342 287 344 289
rect 346 287 348 289
rect 342 285 348 287
rect 561 289 567 291
rect 561 287 563 289
rect 565 287 567 289
rect 561 285 567 287
rect 609 289 615 291
rect 609 287 611 289
rect 613 287 615 289
rect 609 285 615 287
rect 828 289 834 291
rect 828 287 830 289
rect 832 287 834 289
rect 828 285 834 287
rect 35 157 41 159
rect 35 155 37 157
rect 39 155 41 157
rect 35 153 41 155
rect 75 157 81 159
rect 75 155 77 157
rect 79 155 81 157
rect 75 153 81 155
rect 294 157 300 159
rect 294 155 296 157
rect 298 155 300 157
rect 294 153 300 155
rect 342 157 348 159
rect 342 155 344 157
rect 346 155 348 157
rect 342 153 348 155
rect 561 157 567 159
rect 561 155 563 157
rect 565 155 567 157
rect 561 153 567 155
rect 609 157 615 159
rect 609 155 611 157
rect 613 155 615 157
rect 609 153 615 155
rect 828 157 834 159
rect 828 155 830 157
rect 832 155 834 157
rect 828 153 834 155
rect 35 145 41 147
rect 35 143 37 145
rect 39 143 41 145
rect 35 141 41 143
rect 75 145 81 147
rect 75 143 77 145
rect 79 143 81 145
rect 75 141 81 143
rect 294 145 300 147
rect 294 143 296 145
rect 298 143 300 145
rect 294 141 300 143
rect 342 145 348 147
rect 342 143 344 145
rect 346 143 348 145
rect 342 141 348 143
rect 561 145 567 147
rect 561 143 563 145
rect 565 143 567 145
rect 561 141 567 143
rect 609 145 615 147
rect 609 143 611 145
rect 613 143 615 145
rect 609 141 615 143
rect 828 145 834 147
rect 828 143 830 145
rect 832 143 834 145
rect 828 141 834 143
rect 35 13 41 15
rect 35 11 37 13
rect 39 11 41 13
rect 35 9 41 11
rect 75 13 81 15
rect 75 11 77 13
rect 79 11 81 13
rect 75 9 81 11
rect 294 13 300 15
rect 294 11 296 13
rect 298 11 300 13
rect 294 9 300 11
rect 342 13 348 15
rect 342 11 344 13
rect 346 11 348 13
rect 342 9 348 11
rect 561 13 567 15
rect 561 11 563 13
rect 565 11 567 13
rect 561 9 567 11
rect 609 13 615 15
rect 609 11 611 13
rect 613 11 615 13
rect 609 9 615 11
rect 828 13 834 15
rect 828 11 830 13
rect 832 11 834 13
rect 828 9 834 11
rect 458 1 464 3
rect 458 -1 460 1
rect 462 -1 464 1
rect 458 -3 464 -1
rect 696 1 702 3
rect 696 -1 698 1
rect 700 -1 702 1
rect 696 -3 702 -1
rect 458 -131 464 -129
rect 458 -133 460 -131
rect 462 -133 464 -131
rect 458 -135 464 -133
rect 696 -131 702 -129
rect 696 -133 698 -131
rect 700 -133 702 -131
rect 696 -135 702 -133
rect 458 -143 464 -141
rect 458 -145 460 -143
rect 462 -145 464 -143
rect 458 -147 464 -145
rect 696 -143 702 -141
rect 696 -145 698 -143
rect 700 -145 702 -143
rect 696 -147 702 -145
rect 458 -275 464 -273
rect 458 -277 460 -275
rect 462 -277 464 -275
rect 458 -279 464 -277
rect 696 -275 702 -273
rect 696 -277 698 -275
rect 700 -277 702 -275
rect 696 -279 702 -277
<< nmos >>
rect 13 235 15 246
rect 20 235 22 246
rect 33 237 35 246
rect 53 235 55 246
rect 60 235 62 246
rect 73 237 75 246
rect 93 228 95 241
rect 103 231 105 241
rect 113 234 115 248
rect 123 234 125 248
rect 143 228 145 248
rect 150 228 152 248
rect 161 228 163 242
rect 183 228 185 242
rect 194 228 196 248
rect 201 228 203 248
rect 221 234 223 248
rect 231 234 233 248
rect 272 242 274 248
rect 282 242 284 248
rect 241 231 243 241
rect 251 228 253 241
rect 292 239 294 248
rect 320 235 322 246
rect 327 235 329 246
rect 340 237 342 246
rect 360 228 362 241
rect 370 231 372 241
rect 380 234 382 248
rect 390 234 392 248
rect 410 228 412 248
rect 417 228 419 248
rect 428 228 430 242
rect 450 228 452 242
rect 461 228 463 248
rect 468 228 470 248
rect 488 234 490 248
rect 498 234 500 248
rect 539 242 541 248
rect 549 242 551 248
rect 508 231 510 241
rect 518 228 520 241
rect 559 239 561 248
rect 587 235 589 246
rect 594 235 596 246
rect 607 237 609 246
rect 627 228 629 241
rect 637 231 639 241
rect 647 234 649 248
rect 657 234 659 248
rect 677 228 679 248
rect 684 228 686 248
rect 695 228 697 242
rect 717 228 719 242
rect 728 228 730 248
rect 735 228 737 248
rect 755 234 757 248
rect 765 234 767 248
rect 806 242 808 248
rect 816 242 818 248
rect 775 231 777 241
rect 785 228 787 241
rect 826 239 828 248
rect 13 198 15 209
rect 20 198 22 209
rect 33 198 35 207
rect 53 198 55 209
rect 60 198 62 209
rect 73 198 75 207
rect 93 203 95 216
rect 103 203 105 213
rect 113 196 115 210
rect 123 196 125 210
rect 143 196 145 216
rect 150 196 152 216
rect 161 202 163 216
rect 183 202 185 216
rect 194 196 196 216
rect 201 196 203 216
rect 221 196 223 210
rect 231 196 233 210
rect 241 203 243 213
rect 251 203 253 216
rect 272 196 274 202
rect 282 196 284 202
rect 292 196 294 205
rect 320 198 322 209
rect 327 198 329 209
rect 340 198 342 207
rect 360 203 362 216
rect 370 203 372 213
rect 380 196 382 210
rect 390 196 392 210
rect 410 196 412 216
rect 417 196 419 216
rect 428 202 430 216
rect 450 202 452 216
rect 461 196 463 216
rect 468 196 470 216
rect 488 196 490 210
rect 498 196 500 210
rect 508 203 510 213
rect 518 203 520 216
rect 539 196 541 202
rect 549 196 551 202
rect 559 196 561 205
rect 587 198 589 209
rect 594 198 596 209
rect 607 198 609 207
rect 627 203 629 216
rect 637 203 639 213
rect 647 196 649 210
rect 657 196 659 210
rect 677 196 679 216
rect 684 196 686 216
rect 695 202 697 216
rect 717 202 719 216
rect 728 196 730 216
rect 735 196 737 216
rect 755 196 757 210
rect 765 196 767 210
rect 775 203 777 213
rect 785 203 787 216
rect 806 196 808 202
rect 816 196 818 202
rect 826 196 828 205
rect 13 91 15 102
rect 20 91 22 102
rect 33 93 35 102
rect 53 91 55 102
rect 60 91 62 102
rect 73 93 75 102
rect 93 84 95 97
rect 103 87 105 97
rect 113 90 115 104
rect 123 90 125 104
rect 143 84 145 104
rect 150 84 152 104
rect 161 84 163 98
rect 183 84 185 98
rect 194 84 196 104
rect 201 84 203 104
rect 221 90 223 104
rect 231 90 233 104
rect 272 98 274 104
rect 282 98 284 104
rect 241 87 243 97
rect 251 84 253 97
rect 292 95 294 104
rect 320 91 322 102
rect 327 91 329 102
rect 340 93 342 102
rect 360 84 362 97
rect 370 87 372 97
rect 380 90 382 104
rect 390 90 392 104
rect 410 84 412 104
rect 417 84 419 104
rect 428 84 430 98
rect 450 84 452 98
rect 461 84 463 104
rect 468 84 470 104
rect 488 90 490 104
rect 498 90 500 104
rect 539 98 541 104
rect 549 98 551 104
rect 508 87 510 97
rect 518 84 520 97
rect 559 95 561 104
rect 587 91 589 102
rect 594 91 596 102
rect 607 93 609 102
rect 627 84 629 97
rect 637 87 639 97
rect 647 90 649 104
rect 657 90 659 104
rect 677 84 679 104
rect 684 84 686 104
rect 695 84 697 98
rect 717 84 719 98
rect 728 84 730 104
rect 735 84 737 104
rect 755 90 757 104
rect 765 90 767 104
rect 806 98 808 104
rect 816 98 818 104
rect 775 87 777 97
rect 785 84 787 97
rect 826 95 828 104
rect 13 54 15 65
rect 20 54 22 65
rect 33 54 35 63
rect 53 54 55 65
rect 60 54 62 65
rect 73 54 75 63
rect 93 59 95 72
rect 103 59 105 69
rect 113 52 115 66
rect 123 52 125 66
rect 143 52 145 72
rect 150 52 152 72
rect 161 58 163 72
rect 183 58 185 72
rect 194 52 196 72
rect 201 52 203 72
rect 221 52 223 66
rect 231 52 233 66
rect 241 59 243 69
rect 251 59 253 72
rect 272 52 274 58
rect 282 52 284 58
rect 292 52 294 61
rect 320 54 322 65
rect 327 54 329 65
rect 340 54 342 63
rect 360 59 362 72
rect 370 59 372 69
rect 380 52 382 66
rect 390 52 392 66
rect 410 52 412 72
rect 417 52 419 72
rect 428 58 430 72
rect 450 58 452 72
rect 461 52 463 72
rect 468 52 470 72
rect 488 52 490 66
rect 498 52 500 66
rect 508 59 510 69
rect 518 59 520 72
rect 539 52 541 58
rect 549 52 551 58
rect 559 52 561 61
rect 587 54 589 65
rect 594 54 596 65
rect 607 54 609 63
rect 627 59 629 72
rect 637 59 639 69
rect 647 52 649 66
rect 657 52 659 66
rect 677 52 679 72
rect 684 52 686 72
rect 695 58 697 72
rect 717 58 719 72
rect 728 52 730 72
rect 735 52 737 72
rect 755 52 757 66
rect 765 52 767 66
rect 775 59 777 69
rect 785 59 787 72
rect 806 52 808 58
rect 816 52 818 58
rect 826 52 828 61
rect 431 -49 433 -40
rect 447 -54 449 -45
rect 457 -54 459 -45
rect 467 -57 469 -45
rect 474 -57 476 -45
rect 495 -60 497 -47
rect 505 -57 507 -47
rect 515 -54 517 -40
rect 525 -54 527 -40
rect 545 -60 547 -40
rect 552 -60 554 -40
rect 563 -60 565 -46
rect 585 -60 587 -46
rect 596 -60 598 -40
rect 603 -60 605 -40
rect 623 -54 625 -40
rect 633 -54 635 -40
rect 674 -46 676 -40
rect 684 -46 686 -40
rect 643 -57 645 -47
rect 653 -60 655 -47
rect 694 -49 696 -40
rect 717 -52 719 -46
rect 727 -54 729 -46
rect 734 -54 736 -46
rect 744 -54 746 -46
rect 751 -54 753 -46
rect 761 -54 763 -45
rect 781 -52 783 -46
rect 791 -54 793 -46
rect 798 -54 800 -46
rect 808 -54 810 -46
rect 815 -54 817 -46
rect 825 -54 827 -45
rect 431 -92 433 -83
rect 447 -87 449 -78
rect 457 -87 459 -78
rect 467 -87 469 -75
rect 474 -87 476 -75
rect 495 -85 497 -72
rect 505 -85 507 -75
rect 515 -92 517 -78
rect 525 -92 527 -78
rect 545 -92 547 -72
rect 552 -92 554 -72
rect 563 -86 565 -72
rect 585 -86 587 -72
rect 596 -92 598 -72
rect 603 -92 605 -72
rect 623 -92 625 -78
rect 633 -92 635 -78
rect 643 -85 645 -75
rect 653 -85 655 -72
rect 674 -92 676 -86
rect 684 -92 686 -86
rect 694 -92 696 -83
rect 717 -86 719 -80
rect 727 -86 729 -78
rect 734 -86 736 -78
rect 744 -86 746 -78
rect 751 -86 753 -78
rect 761 -87 763 -78
rect 781 -86 783 -80
rect 791 -86 793 -78
rect 798 -86 800 -78
rect 808 -86 810 -78
rect 815 -86 817 -78
rect 825 -87 827 -78
rect 431 -193 433 -184
rect 447 -198 449 -189
rect 457 -198 459 -189
rect 467 -201 469 -189
rect 474 -201 476 -189
rect 495 -204 497 -191
rect 505 -201 507 -191
rect 515 -198 517 -184
rect 525 -198 527 -184
rect 545 -204 547 -184
rect 552 -204 554 -184
rect 563 -204 565 -190
rect 585 -204 587 -190
rect 596 -204 598 -184
rect 603 -204 605 -184
rect 623 -198 625 -184
rect 633 -198 635 -184
rect 674 -190 676 -184
rect 684 -190 686 -184
rect 643 -201 645 -191
rect 653 -204 655 -191
rect 694 -193 696 -184
rect 717 -196 719 -190
rect 727 -198 729 -190
rect 734 -198 736 -190
rect 744 -198 746 -190
rect 751 -198 753 -190
rect 761 -198 763 -189
rect 781 -196 783 -190
rect 791 -198 793 -190
rect 798 -198 800 -190
rect 808 -198 810 -190
rect 815 -198 817 -190
rect 825 -198 827 -189
rect 431 -236 433 -227
rect 447 -231 449 -222
rect 457 -231 459 -222
rect 467 -231 469 -219
rect 474 -231 476 -219
rect 495 -229 497 -216
rect 505 -229 507 -219
rect 515 -236 517 -222
rect 525 -236 527 -222
rect 545 -236 547 -216
rect 552 -236 554 -216
rect 563 -230 565 -216
rect 585 -230 587 -216
rect 596 -236 598 -216
rect 603 -236 605 -216
rect 623 -236 625 -222
rect 633 -236 635 -222
rect 643 -229 645 -219
rect 653 -229 655 -216
rect 674 -236 676 -230
rect 684 -236 686 -230
rect 694 -236 696 -227
rect 717 -230 719 -224
rect 727 -230 729 -222
rect 734 -230 736 -222
rect 744 -230 746 -222
rect 751 -230 753 -222
rect 761 -231 763 -222
rect 781 -230 783 -224
rect 791 -230 793 -222
rect 798 -230 800 -222
rect 808 -230 810 -222
rect 815 -230 817 -222
rect 825 -231 827 -222
<< pmos >>
rect 13 268 15 281
rect 23 268 25 281
rect 33 261 35 279
rect 53 268 55 281
rect 63 268 65 281
rect 73 261 75 279
rect 93 263 95 288
rect 106 263 108 276
rect 116 260 118 285
rect 123 260 125 285
rect 141 260 143 288
rect 151 260 153 288
rect 161 260 163 288
rect 183 260 185 288
rect 193 260 195 288
rect 203 260 205 288
rect 221 260 223 285
rect 228 260 230 285
rect 238 263 240 276
rect 251 263 253 288
rect 272 267 274 288
rect 279 267 281 288
rect 292 260 294 278
rect 320 268 322 281
rect 330 268 332 281
rect 340 261 342 279
rect 360 263 362 288
rect 373 263 375 276
rect 383 260 385 285
rect 390 260 392 285
rect 408 260 410 288
rect 418 260 420 288
rect 428 260 430 288
rect 450 260 452 288
rect 460 260 462 288
rect 470 260 472 288
rect 488 260 490 285
rect 495 260 497 285
rect 505 263 507 276
rect 518 263 520 288
rect 539 267 541 288
rect 546 267 548 288
rect 559 260 561 278
rect 587 268 589 281
rect 597 268 599 281
rect 607 261 609 279
rect 627 263 629 288
rect 640 263 642 276
rect 650 260 652 285
rect 657 260 659 285
rect 675 260 677 288
rect 685 260 687 288
rect 695 260 697 288
rect 717 260 719 288
rect 727 260 729 288
rect 737 260 739 288
rect 755 260 757 285
rect 762 260 764 285
rect 772 263 774 276
rect 785 263 787 288
rect 806 267 808 288
rect 813 267 815 288
rect 826 260 828 278
rect 13 163 15 176
rect 23 163 25 176
rect 33 165 35 183
rect 53 163 55 176
rect 63 163 65 176
rect 73 165 75 183
rect 93 156 95 181
rect 106 168 108 181
rect 116 159 118 184
rect 123 159 125 184
rect 141 156 143 184
rect 151 156 153 184
rect 161 156 163 184
rect 183 156 185 184
rect 193 156 195 184
rect 203 156 205 184
rect 221 159 223 184
rect 228 159 230 184
rect 238 168 240 181
rect 251 156 253 181
rect 272 156 274 177
rect 279 156 281 177
rect 292 166 294 184
rect 320 163 322 176
rect 330 163 332 176
rect 340 165 342 183
rect 360 156 362 181
rect 373 168 375 181
rect 383 159 385 184
rect 390 159 392 184
rect 408 156 410 184
rect 418 156 420 184
rect 428 156 430 184
rect 450 156 452 184
rect 460 156 462 184
rect 470 156 472 184
rect 488 159 490 184
rect 495 159 497 184
rect 505 168 507 181
rect 518 156 520 181
rect 539 156 541 177
rect 546 156 548 177
rect 559 166 561 184
rect 587 163 589 176
rect 597 163 599 176
rect 607 165 609 183
rect 627 156 629 181
rect 640 168 642 181
rect 650 159 652 184
rect 657 159 659 184
rect 675 156 677 184
rect 685 156 687 184
rect 695 156 697 184
rect 717 156 719 184
rect 727 156 729 184
rect 737 156 739 184
rect 755 159 757 184
rect 762 159 764 184
rect 772 168 774 181
rect 785 156 787 181
rect 806 156 808 177
rect 813 156 815 177
rect 826 166 828 184
rect 13 124 15 137
rect 23 124 25 137
rect 33 117 35 135
rect 53 124 55 137
rect 63 124 65 137
rect 73 117 75 135
rect 93 119 95 144
rect 106 119 108 132
rect 116 116 118 141
rect 123 116 125 141
rect 141 116 143 144
rect 151 116 153 144
rect 161 116 163 144
rect 183 116 185 144
rect 193 116 195 144
rect 203 116 205 144
rect 221 116 223 141
rect 228 116 230 141
rect 238 119 240 132
rect 251 119 253 144
rect 272 123 274 144
rect 279 123 281 144
rect 292 116 294 134
rect 320 124 322 137
rect 330 124 332 137
rect 340 117 342 135
rect 360 119 362 144
rect 373 119 375 132
rect 383 116 385 141
rect 390 116 392 141
rect 408 116 410 144
rect 418 116 420 144
rect 428 116 430 144
rect 450 116 452 144
rect 460 116 462 144
rect 470 116 472 144
rect 488 116 490 141
rect 495 116 497 141
rect 505 119 507 132
rect 518 119 520 144
rect 539 123 541 144
rect 546 123 548 144
rect 559 116 561 134
rect 587 124 589 137
rect 597 124 599 137
rect 607 117 609 135
rect 627 119 629 144
rect 640 119 642 132
rect 650 116 652 141
rect 657 116 659 141
rect 675 116 677 144
rect 685 116 687 144
rect 695 116 697 144
rect 717 116 719 144
rect 727 116 729 144
rect 737 116 739 144
rect 755 116 757 141
rect 762 116 764 141
rect 772 119 774 132
rect 785 119 787 144
rect 806 123 808 144
rect 813 123 815 144
rect 826 116 828 134
rect 13 19 15 32
rect 23 19 25 32
rect 33 21 35 39
rect 53 19 55 32
rect 63 19 65 32
rect 73 21 75 39
rect 93 12 95 37
rect 106 24 108 37
rect 116 15 118 40
rect 123 15 125 40
rect 141 12 143 40
rect 151 12 153 40
rect 161 12 163 40
rect 183 12 185 40
rect 193 12 195 40
rect 203 12 205 40
rect 221 15 223 40
rect 228 15 230 40
rect 238 24 240 37
rect 251 12 253 37
rect 272 12 274 33
rect 279 12 281 33
rect 292 22 294 40
rect 320 19 322 32
rect 330 19 332 32
rect 340 21 342 39
rect 360 12 362 37
rect 373 24 375 37
rect 383 15 385 40
rect 390 15 392 40
rect 408 12 410 40
rect 418 12 420 40
rect 428 12 430 40
rect 450 12 452 40
rect 460 12 462 40
rect 470 12 472 40
rect 488 15 490 40
rect 495 15 497 40
rect 505 24 507 37
rect 518 12 520 37
rect 539 12 541 33
rect 546 12 548 33
rect 559 22 561 40
rect 587 19 589 32
rect 597 19 599 32
rect 607 21 609 39
rect 627 12 629 37
rect 640 24 642 37
rect 650 15 652 40
rect 657 15 659 40
rect 675 12 677 40
rect 685 12 687 40
rect 695 12 697 40
rect 717 12 719 40
rect 727 12 729 40
rect 737 12 739 40
rect 755 15 757 40
rect 762 15 764 40
rect 772 24 774 37
rect 785 12 787 37
rect 806 12 808 33
rect 813 12 815 33
rect 826 22 828 40
rect 439 -27 441 0
rect 455 -27 457 -9
rect 465 -27 467 -9
rect 475 -27 477 0
rect 495 -25 497 0
rect 508 -25 510 -12
rect 518 -28 520 -3
rect 525 -28 527 -3
rect 543 -28 545 0
rect 553 -28 555 0
rect 563 -28 565 0
rect 585 -28 587 0
rect 595 -28 597 0
rect 605 -28 607 0
rect 623 -28 625 -3
rect 630 -28 632 -3
rect 640 -25 642 -12
rect 653 -25 655 0
rect 674 -21 676 0
rect 681 -21 683 0
rect 694 -28 696 -10
rect 727 -16 729 0
rect 734 -16 736 0
rect 744 -16 746 0
rect 751 -16 753 0
rect 717 -28 719 -20
rect 761 -18 763 0
rect 791 -16 793 0
rect 798 -16 800 0
rect 808 -16 810 0
rect 815 -16 817 0
rect 781 -28 783 -20
rect 825 -18 827 0
rect 439 -132 441 -105
rect 455 -123 457 -105
rect 465 -123 467 -105
rect 475 -132 477 -105
rect 495 -132 497 -107
rect 508 -120 510 -107
rect 518 -129 520 -104
rect 525 -129 527 -104
rect 543 -132 545 -104
rect 553 -132 555 -104
rect 563 -132 565 -104
rect 585 -132 587 -104
rect 595 -132 597 -104
rect 605 -132 607 -104
rect 623 -129 625 -104
rect 630 -129 632 -104
rect 640 -120 642 -107
rect 653 -132 655 -107
rect 674 -132 676 -111
rect 681 -132 683 -111
rect 694 -122 696 -104
rect 717 -112 719 -104
rect 781 -112 783 -104
rect 727 -132 729 -116
rect 734 -132 736 -116
rect 744 -132 746 -116
rect 751 -132 753 -116
rect 761 -132 763 -114
rect 791 -132 793 -116
rect 798 -132 800 -116
rect 808 -132 810 -116
rect 815 -132 817 -116
rect 825 -132 827 -114
rect 439 -171 441 -144
rect 455 -171 457 -153
rect 465 -171 467 -153
rect 475 -171 477 -144
rect 495 -169 497 -144
rect 508 -169 510 -156
rect 518 -172 520 -147
rect 525 -172 527 -147
rect 543 -172 545 -144
rect 553 -172 555 -144
rect 563 -172 565 -144
rect 585 -172 587 -144
rect 595 -172 597 -144
rect 605 -172 607 -144
rect 623 -172 625 -147
rect 630 -172 632 -147
rect 640 -169 642 -156
rect 653 -169 655 -144
rect 674 -165 676 -144
rect 681 -165 683 -144
rect 694 -172 696 -154
rect 727 -160 729 -144
rect 734 -160 736 -144
rect 744 -160 746 -144
rect 751 -160 753 -144
rect 717 -172 719 -164
rect 761 -162 763 -144
rect 791 -160 793 -144
rect 798 -160 800 -144
rect 808 -160 810 -144
rect 815 -160 817 -144
rect 781 -172 783 -164
rect 825 -162 827 -144
rect 439 -276 441 -249
rect 455 -267 457 -249
rect 465 -267 467 -249
rect 475 -276 477 -249
rect 495 -276 497 -251
rect 508 -264 510 -251
rect 518 -273 520 -248
rect 525 -273 527 -248
rect 543 -276 545 -248
rect 553 -276 555 -248
rect 563 -276 565 -248
rect 585 -276 587 -248
rect 595 -276 597 -248
rect 605 -276 607 -248
rect 623 -273 625 -248
rect 630 -273 632 -248
rect 640 -264 642 -251
rect 653 -276 655 -251
rect 674 -276 676 -255
rect 681 -276 683 -255
rect 694 -266 696 -248
rect 717 -256 719 -248
rect 781 -256 783 -248
rect 727 -276 729 -260
rect 734 -276 736 -260
rect 744 -276 746 -260
rect 751 -276 753 -260
rect 761 -276 763 -258
rect 791 -276 793 -260
rect 798 -276 800 -260
rect 808 -276 810 -260
rect 815 -276 817 -260
rect 825 -276 827 -258
<< polyct0 >>
rect 31 253 33 255
rect 71 253 73 255
rect 101 256 103 258
rect 95 246 97 248
rect 151 253 153 255
rect 161 253 163 255
rect 183 253 185 255
rect 193 253 195 255
rect 243 256 245 258
rect 290 253 292 255
rect 249 246 251 248
rect 338 253 340 255
rect 368 256 370 258
rect 362 246 364 248
rect 418 253 420 255
rect 428 253 430 255
rect 450 253 452 255
rect 460 253 462 255
rect 510 256 512 258
rect 557 253 559 255
rect 516 246 518 248
rect 605 253 607 255
rect 635 256 637 258
rect 629 246 631 248
rect 685 253 687 255
rect 695 253 697 255
rect 717 253 719 255
rect 727 253 729 255
rect 777 256 779 258
rect 824 253 826 255
rect 783 246 785 248
rect 31 189 33 191
rect 71 189 73 191
rect 95 196 97 198
rect 101 186 103 188
rect 151 189 153 191
rect 161 189 163 191
rect 183 189 185 191
rect 193 189 195 191
rect 249 196 251 198
rect 243 186 245 188
rect 290 189 292 191
rect 338 189 340 191
rect 362 196 364 198
rect 368 186 370 188
rect 418 189 420 191
rect 428 189 430 191
rect 450 189 452 191
rect 460 189 462 191
rect 516 196 518 198
rect 510 186 512 188
rect 557 189 559 191
rect 605 189 607 191
rect 629 196 631 198
rect 635 186 637 188
rect 685 189 687 191
rect 695 189 697 191
rect 717 189 719 191
rect 727 189 729 191
rect 783 196 785 198
rect 777 186 779 188
rect 824 189 826 191
rect 31 109 33 111
rect 71 109 73 111
rect 101 112 103 114
rect 95 102 97 104
rect 151 109 153 111
rect 161 109 163 111
rect 183 109 185 111
rect 193 109 195 111
rect 243 112 245 114
rect 290 109 292 111
rect 249 102 251 104
rect 338 109 340 111
rect 368 112 370 114
rect 362 102 364 104
rect 418 109 420 111
rect 428 109 430 111
rect 450 109 452 111
rect 460 109 462 111
rect 510 112 512 114
rect 557 109 559 111
rect 516 102 518 104
rect 605 109 607 111
rect 635 112 637 114
rect 629 102 631 104
rect 685 109 687 111
rect 695 109 697 111
rect 717 109 719 111
rect 727 109 729 111
rect 777 112 779 114
rect 824 109 826 111
rect 783 102 785 104
rect 31 45 33 47
rect 71 45 73 47
rect 95 52 97 54
rect 101 42 103 44
rect 151 45 153 47
rect 161 45 163 47
rect 183 45 185 47
rect 193 45 195 47
rect 249 52 251 54
rect 243 42 245 44
rect 290 45 292 47
rect 338 45 340 47
rect 362 52 364 54
rect 368 42 370 44
rect 418 45 420 47
rect 428 45 430 47
rect 450 45 452 47
rect 460 45 462 47
rect 516 52 518 54
rect 510 42 512 44
rect 557 45 559 47
rect 605 45 607 47
rect 629 52 631 54
rect 635 42 637 44
rect 685 45 687 47
rect 695 45 697 47
rect 717 45 719 47
rect 727 45 729 47
rect 783 52 785 54
rect 777 42 779 44
rect 824 45 826 47
rect 463 -35 465 -33
rect 473 -34 475 -32
rect 503 -32 505 -30
rect 497 -42 499 -40
rect 553 -35 555 -33
rect 563 -35 565 -33
rect 585 -35 587 -33
rect 595 -35 597 -33
rect 645 -32 647 -30
rect 692 -35 694 -33
rect 651 -42 653 -40
rect 735 -25 737 -23
rect 742 -41 744 -39
rect 760 -40 762 -38
rect 799 -25 801 -23
rect 806 -41 808 -39
rect 824 -40 826 -38
rect 497 -92 499 -90
rect 463 -99 465 -97
rect 473 -100 475 -98
rect 503 -102 505 -100
rect 553 -99 555 -97
rect 563 -99 565 -97
rect 585 -99 587 -97
rect 595 -99 597 -97
rect 651 -92 653 -90
rect 645 -102 647 -100
rect 692 -99 694 -97
rect 742 -93 744 -91
rect 760 -94 762 -92
rect 735 -109 737 -107
rect 806 -93 808 -91
rect 824 -94 826 -92
rect 799 -109 801 -107
rect 463 -179 465 -177
rect 473 -178 475 -176
rect 503 -176 505 -174
rect 497 -186 499 -184
rect 553 -179 555 -177
rect 563 -179 565 -177
rect 585 -179 587 -177
rect 595 -179 597 -177
rect 645 -176 647 -174
rect 692 -179 694 -177
rect 651 -186 653 -184
rect 735 -169 737 -167
rect 742 -185 744 -183
rect 760 -184 762 -182
rect 799 -169 801 -167
rect 806 -185 808 -183
rect 824 -184 826 -182
rect 497 -236 499 -234
rect 463 -243 465 -241
rect 473 -244 475 -242
rect 503 -246 505 -244
rect 553 -243 555 -241
rect 563 -243 565 -241
rect 585 -243 587 -241
rect 595 -243 597 -241
rect 651 -236 653 -234
rect 645 -246 647 -244
rect 692 -243 694 -241
rect 742 -237 744 -235
rect 760 -238 762 -236
rect 735 -253 737 -251
rect 806 -237 808 -235
rect 824 -238 826 -236
rect 799 -253 801 -251
<< polyct1 >>
rect 11 261 13 263
rect 51 261 53 263
rect 21 253 23 255
rect 61 253 63 255
rect 115 253 117 255
rect 134 253 136 255
rect 141 253 143 255
rect 203 253 205 255
rect 210 253 212 255
rect 229 253 231 255
rect 270 260 272 262
rect 318 261 320 263
rect 280 253 282 255
rect 328 253 330 255
rect 382 253 384 255
rect 401 253 403 255
rect 408 253 410 255
rect 470 253 472 255
rect 477 253 479 255
rect 496 253 498 255
rect 537 260 539 262
rect 585 261 587 263
rect 547 253 549 255
rect 595 253 597 255
rect 649 253 651 255
rect 668 253 670 255
rect 675 253 677 255
rect 737 253 739 255
rect 744 253 746 255
rect 763 253 765 255
rect 804 260 806 262
rect 814 253 816 255
rect 21 189 23 191
rect 11 181 13 183
rect 61 189 63 191
rect 51 181 53 183
rect 115 189 117 191
rect 134 189 136 191
rect 141 189 143 191
rect 203 189 205 191
rect 210 189 212 191
rect 229 189 231 191
rect 280 189 282 191
rect 270 182 272 184
rect 328 189 330 191
rect 318 181 320 183
rect 382 189 384 191
rect 401 189 403 191
rect 408 189 410 191
rect 470 189 472 191
rect 477 189 479 191
rect 496 189 498 191
rect 547 189 549 191
rect 537 182 539 184
rect 595 189 597 191
rect 585 181 587 183
rect 649 189 651 191
rect 668 189 670 191
rect 675 189 677 191
rect 737 189 739 191
rect 744 189 746 191
rect 763 189 765 191
rect 814 189 816 191
rect 804 182 806 184
rect 11 117 13 119
rect 51 117 53 119
rect 21 109 23 111
rect 61 109 63 111
rect 115 109 117 111
rect 134 109 136 111
rect 141 109 143 111
rect 203 109 205 111
rect 210 109 212 111
rect 229 109 231 111
rect 270 116 272 118
rect 318 117 320 119
rect 280 109 282 111
rect 328 109 330 111
rect 382 109 384 111
rect 401 109 403 111
rect 408 109 410 111
rect 470 109 472 111
rect 477 109 479 111
rect 496 109 498 111
rect 537 116 539 118
rect 585 117 587 119
rect 547 109 549 111
rect 595 109 597 111
rect 649 109 651 111
rect 668 109 670 111
rect 675 109 677 111
rect 737 109 739 111
rect 744 109 746 111
rect 763 109 765 111
rect 804 116 806 118
rect 814 109 816 111
rect 21 45 23 47
rect 11 37 13 39
rect 61 45 63 47
rect 51 37 53 39
rect 115 45 117 47
rect 134 45 136 47
rect 141 45 143 47
rect 203 45 205 47
rect 210 45 212 47
rect 229 45 231 47
rect 280 45 282 47
rect 270 38 272 40
rect 328 45 330 47
rect 318 37 320 39
rect 382 45 384 47
rect 401 45 403 47
rect 408 45 410 47
rect 470 45 472 47
rect 477 45 479 47
rect 496 45 498 47
rect 547 45 549 47
rect 537 38 539 40
rect 595 45 597 47
rect 585 37 587 39
rect 649 45 651 47
rect 668 45 670 47
rect 675 45 677 47
rect 737 45 739 47
rect 744 45 746 47
rect 763 45 765 47
rect 814 45 816 47
rect 804 38 806 40
rect 426 -27 428 -25
rect 442 -40 444 -38
rect 517 -35 519 -33
rect 536 -35 538 -33
rect 543 -35 545 -33
rect 605 -35 607 -33
rect 612 -35 614 -33
rect 631 -35 633 -33
rect 672 -28 674 -26
rect 712 -15 714 -13
rect 682 -35 684 -33
rect 776 -15 778 -13
rect 725 -35 727 -33
rect 752 -30 754 -28
rect 789 -35 791 -33
rect 816 -30 818 -28
rect 442 -94 444 -92
rect 426 -107 428 -105
rect 517 -99 519 -97
rect 536 -99 538 -97
rect 543 -99 545 -97
rect 605 -99 607 -97
rect 612 -99 614 -97
rect 631 -99 633 -97
rect 682 -99 684 -97
rect 672 -106 674 -104
rect 725 -99 727 -97
rect 752 -104 754 -102
rect 789 -99 791 -97
rect 712 -119 714 -117
rect 816 -104 818 -102
rect 776 -119 778 -117
rect 426 -171 428 -169
rect 442 -184 444 -182
rect 517 -179 519 -177
rect 536 -179 538 -177
rect 543 -179 545 -177
rect 605 -179 607 -177
rect 612 -179 614 -177
rect 631 -179 633 -177
rect 672 -172 674 -170
rect 712 -159 714 -157
rect 682 -179 684 -177
rect 776 -159 778 -157
rect 725 -179 727 -177
rect 752 -174 754 -172
rect 789 -179 791 -177
rect 816 -174 818 -172
rect 442 -238 444 -236
rect 426 -251 428 -249
rect 517 -243 519 -241
rect 536 -243 538 -241
rect 543 -243 545 -241
rect 605 -243 607 -241
rect 612 -243 614 -241
rect 631 -243 633 -241
rect 682 -243 684 -241
rect 672 -250 674 -248
rect 725 -243 727 -241
rect 752 -248 754 -246
rect 789 -243 791 -241
rect 712 -263 714 -261
rect 816 -248 818 -246
rect 776 -263 778 -261
<< ndifct0 >>
rect 8 237 10 239
rect 48 237 50 239
rect 98 233 100 235
rect 108 236 110 238
rect 118 244 120 246
rect 128 244 130 246
rect 128 237 130 239
rect 138 237 140 239
rect 155 230 157 232
rect 189 230 191 232
rect 216 244 218 246
rect 206 237 208 239
rect 216 237 218 239
rect 226 244 228 246
rect 277 244 279 246
rect 236 236 238 238
rect 246 233 248 235
rect 267 231 269 233
rect 315 237 317 239
rect 286 231 288 233
rect 365 233 367 235
rect 375 236 377 238
rect 385 244 387 246
rect 395 244 397 246
rect 395 237 397 239
rect 405 237 407 239
rect 422 230 424 232
rect 456 230 458 232
rect 483 244 485 246
rect 473 237 475 239
rect 483 237 485 239
rect 493 244 495 246
rect 544 244 546 246
rect 503 236 505 238
rect 513 233 515 235
rect 534 231 536 233
rect 582 237 584 239
rect 553 231 555 233
rect 632 233 634 235
rect 642 236 644 238
rect 652 244 654 246
rect 662 244 664 246
rect 662 237 664 239
rect 672 237 674 239
rect 689 230 691 232
rect 723 230 725 232
rect 750 244 752 246
rect 740 237 742 239
rect 750 237 752 239
rect 760 244 762 246
rect 811 244 813 246
rect 770 236 772 238
rect 780 233 782 235
rect 801 231 803 233
rect 820 231 822 233
rect 8 205 10 207
rect 48 205 50 207
rect 98 209 100 211
rect 108 206 110 208
rect 118 198 120 200
rect 128 205 130 207
rect 138 205 140 207
rect 128 198 130 200
rect 155 212 157 214
rect 189 212 191 214
rect 206 205 208 207
rect 216 205 218 207
rect 216 198 218 200
rect 226 198 228 200
rect 236 206 238 208
rect 246 209 248 211
rect 267 211 269 213
rect 286 211 288 213
rect 315 205 317 207
rect 277 198 279 200
rect 365 209 367 211
rect 375 206 377 208
rect 385 198 387 200
rect 395 205 397 207
rect 405 205 407 207
rect 395 198 397 200
rect 422 212 424 214
rect 456 212 458 214
rect 473 205 475 207
rect 483 205 485 207
rect 483 198 485 200
rect 493 198 495 200
rect 503 206 505 208
rect 513 209 515 211
rect 534 211 536 213
rect 553 211 555 213
rect 582 205 584 207
rect 544 198 546 200
rect 632 209 634 211
rect 642 206 644 208
rect 652 198 654 200
rect 662 205 664 207
rect 672 205 674 207
rect 662 198 664 200
rect 689 212 691 214
rect 723 212 725 214
rect 740 205 742 207
rect 750 205 752 207
rect 750 198 752 200
rect 760 198 762 200
rect 770 206 772 208
rect 780 209 782 211
rect 801 211 803 213
rect 820 211 822 213
rect 811 198 813 200
rect 8 93 10 95
rect 48 93 50 95
rect 98 89 100 91
rect 108 92 110 94
rect 118 100 120 102
rect 128 100 130 102
rect 128 93 130 95
rect 138 93 140 95
rect 155 86 157 88
rect 189 86 191 88
rect 216 100 218 102
rect 206 93 208 95
rect 216 93 218 95
rect 226 100 228 102
rect 277 100 279 102
rect 236 92 238 94
rect 246 89 248 91
rect 267 87 269 89
rect 315 93 317 95
rect 286 87 288 89
rect 365 89 367 91
rect 375 92 377 94
rect 385 100 387 102
rect 395 100 397 102
rect 395 93 397 95
rect 405 93 407 95
rect 422 86 424 88
rect 456 86 458 88
rect 483 100 485 102
rect 473 93 475 95
rect 483 93 485 95
rect 493 100 495 102
rect 544 100 546 102
rect 503 92 505 94
rect 513 89 515 91
rect 534 87 536 89
rect 582 93 584 95
rect 553 87 555 89
rect 632 89 634 91
rect 642 92 644 94
rect 652 100 654 102
rect 662 100 664 102
rect 662 93 664 95
rect 672 93 674 95
rect 689 86 691 88
rect 723 86 725 88
rect 750 100 752 102
rect 740 93 742 95
rect 750 93 752 95
rect 760 100 762 102
rect 811 100 813 102
rect 770 92 772 94
rect 780 89 782 91
rect 801 87 803 89
rect 820 87 822 89
rect 8 61 10 63
rect 48 61 50 63
rect 98 65 100 67
rect 108 62 110 64
rect 118 54 120 56
rect 128 61 130 63
rect 138 61 140 63
rect 128 54 130 56
rect 155 68 157 70
rect 189 68 191 70
rect 206 61 208 63
rect 216 61 218 63
rect 216 54 218 56
rect 226 54 228 56
rect 236 62 238 64
rect 246 65 248 67
rect 267 67 269 69
rect 286 67 288 69
rect 315 61 317 63
rect 277 54 279 56
rect 365 65 367 67
rect 375 62 377 64
rect 385 54 387 56
rect 395 61 397 63
rect 405 61 407 63
rect 395 54 397 56
rect 422 68 424 70
rect 456 68 458 70
rect 473 61 475 63
rect 483 61 485 63
rect 483 54 485 56
rect 493 54 495 56
rect 503 62 505 64
rect 513 65 515 67
rect 534 67 536 69
rect 553 67 555 69
rect 582 61 584 63
rect 544 54 546 56
rect 632 65 634 67
rect 642 62 644 64
rect 652 54 654 56
rect 662 61 664 63
rect 672 61 674 63
rect 662 54 664 56
rect 689 68 691 70
rect 723 68 725 70
rect 740 61 742 63
rect 750 61 752 63
rect 750 54 752 56
rect 760 54 762 56
rect 770 62 772 64
rect 780 65 782 67
rect 801 67 803 69
rect 820 67 822 69
rect 811 54 813 56
rect 426 -44 428 -42
rect 440 -52 442 -50
rect 452 -49 454 -47
rect 500 -55 502 -53
rect 510 -52 512 -50
rect 520 -44 522 -42
rect 530 -44 532 -42
rect 530 -51 532 -49
rect 540 -51 542 -49
rect 557 -58 559 -56
rect 591 -58 593 -56
rect 618 -44 620 -42
rect 608 -51 610 -49
rect 618 -51 620 -49
rect 628 -44 630 -42
rect 679 -44 681 -42
rect 638 -52 640 -50
rect 648 -55 650 -53
rect 669 -57 671 -55
rect 712 -50 714 -48
rect 722 -50 724 -48
rect 688 -57 690 -55
rect 739 -52 741 -50
rect 756 -52 758 -50
rect 776 -50 778 -48
rect 786 -50 788 -48
rect 803 -52 805 -50
rect 820 -52 822 -50
rect 440 -82 442 -80
rect 426 -90 428 -88
rect 452 -85 454 -83
rect 500 -79 502 -77
rect 510 -82 512 -80
rect 520 -90 522 -88
rect 530 -83 532 -81
rect 540 -83 542 -81
rect 530 -90 532 -88
rect 557 -76 559 -74
rect 591 -76 593 -74
rect 608 -83 610 -81
rect 618 -83 620 -81
rect 618 -90 620 -88
rect 628 -90 630 -88
rect 638 -82 640 -80
rect 648 -79 650 -77
rect 669 -77 671 -75
rect 688 -77 690 -75
rect 679 -90 681 -88
rect 712 -84 714 -82
rect 722 -84 724 -82
rect 739 -82 741 -80
rect 756 -82 758 -80
rect 776 -84 778 -82
rect 786 -84 788 -82
rect 803 -82 805 -80
rect 820 -82 822 -80
rect 426 -188 428 -186
rect 440 -196 442 -194
rect 452 -193 454 -191
rect 500 -199 502 -197
rect 510 -196 512 -194
rect 520 -188 522 -186
rect 530 -188 532 -186
rect 530 -195 532 -193
rect 540 -195 542 -193
rect 557 -202 559 -200
rect 591 -202 593 -200
rect 618 -188 620 -186
rect 608 -195 610 -193
rect 618 -195 620 -193
rect 628 -188 630 -186
rect 679 -188 681 -186
rect 638 -196 640 -194
rect 648 -199 650 -197
rect 669 -201 671 -199
rect 712 -194 714 -192
rect 722 -194 724 -192
rect 688 -201 690 -199
rect 739 -196 741 -194
rect 756 -196 758 -194
rect 776 -194 778 -192
rect 786 -194 788 -192
rect 803 -196 805 -194
rect 820 -196 822 -194
rect 440 -226 442 -224
rect 426 -234 428 -232
rect 452 -229 454 -227
rect 500 -223 502 -221
rect 510 -226 512 -224
rect 520 -234 522 -232
rect 530 -227 532 -225
rect 540 -227 542 -225
rect 530 -234 532 -232
rect 557 -220 559 -218
rect 591 -220 593 -218
rect 608 -227 610 -225
rect 618 -227 620 -225
rect 618 -234 620 -232
rect 628 -234 630 -232
rect 638 -226 640 -224
rect 648 -223 650 -221
rect 669 -221 671 -219
rect 688 -221 690 -219
rect 679 -234 681 -232
rect 712 -228 714 -226
rect 722 -228 724 -226
rect 739 -226 741 -224
rect 756 -226 758 -224
rect 776 -228 778 -226
rect 786 -228 788 -226
rect 803 -226 805 -224
rect 820 -226 822 -224
<< ndifct1 >>
rect 38 239 40 241
rect 78 239 80 241
rect 88 237 90 239
rect 27 227 29 229
rect 67 227 69 229
rect 166 237 168 239
rect 178 237 180 239
rect 256 237 258 239
rect 297 244 299 246
rect 345 239 347 241
rect 355 237 357 239
rect 334 227 336 229
rect 433 237 435 239
rect 445 237 447 239
rect 523 237 525 239
rect 564 244 566 246
rect 612 239 614 241
rect 622 237 624 239
rect 601 227 603 229
rect 700 237 702 239
rect 712 237 714 239
rect 790 237 792 239
rect 831 244 833 246
rect 27 215 29 217
rect 67 215 69 217
rect 38 203 40 205
rect 78 203 80 205
rect 88 205 90 207
rect 166 205 168 207
rect 178 205 180 207
rect 334 215 336 217
rect 256 205 258 207
rect 297 198 299 200
rect 345 203 347 205
rect 355 205 357 207
rect 433 205 435 207
rect 445 205 447 207
rect 601 215 603 217
rect 523 205 525 207
rect 564 198 566 200
rect 612 203 614 205
rect 622 205 624 207
rect 700 205 702 207
rect 712 205 714 207
rect 790 205 792 207
rect 831 198 833 200
rect 38 95 40 97
rect 78 95 80 97
rect 88 93 90 95
rect 27 83 29 85
rect 67 83 69 85
rect 166 93 168 95
rect 178 93 180 95
rect 256 93 258 95
rect 297 100 299 102
rect 345 95 347 97
rect 355 93 357 95
rect 334 83 336 85
rect 433 93 435 95
rect 445 93 447 95
rect 523 93 525 95
rect 564 100 566 102
rect 612 95 614 97
rect 622 93 624 95
rect 601 83 603 85
rect 700 93 702 95
rect 712 93 714 95
rect 790 93 792 95
rect 831 100 833 102
rect 27 71 29 73
rect 67 71 69 73
rect 38 59 40 61
rect 78 59 80 61
rect 88 61 90 63
rect 166 61 168 63
rect 178 61 180 63
rect 334 71 336 73
rect 256 61 258 63
rect 297 54 299 56
rect 345 59 347 61
rect 355 61 357 63
rect 433 61 435 63
rect 445 61 447 63
rect 601 71 603 73
rect 523 61 525 63
rect 564 54 566 56
rect 612 59 614 61
rect 622 61 624 63
rect 700 61 702 63
rect 712 61 714 63
rect 790 61 792 63
rect 831 54 833 56
rect 462 -51 464 -49
rect 490 -51 492 -49
rect 480 -61 482 -59
rect 568 -51 570 -49
rect 580 -51 582 -49
rect 658 -51 660 -49
rect 699 -44 701 -42
rect 766 -49 768 -47
rect 830 -49 832 -47
rect 480 -73 482 -71
rect 462 -83 464 -81
rect 490 -83 492 -81
rect 568 -83 570 -81
rect 580 -83 582 -81
rect 658 -83 660 -81
rect 699 -90 701 -88
rect 766 -85 768 -83
rect 830 -85 832 -83
rect 462 -195 464 -193
rect 490 -195 492 -193
rect 480 -205 482 -203
rect 568 -195 570 -193
rect 580 -195 582 -193
rect 658 -195 660 -193
rect 699 -188 701 -186
rect 766 -193 768 -191
rect 830 -193 832 -191
rect 480 -217 482 -215
rect 462 -227 464 -225
rect 490 -227 492 -225
rect 568 -227 570 -225
rect 580 -227 582 -225
rect 658 -227 660 -225
rect 699 -234 701 -232
rect 766 -229 768 -227
rect 830 -229 832 -227
<< ntiect1 >>
rect 37 287 39 289
rect 77 287 79 289
rect 296 287 298 289
rect 344 287 346 289
rect 563 287 565 289
rect 611 287 613 289
rect 830 287 832 289
rect 37 155 39 157
rect 77 155 79 157
rect 296 155 298 157
rect 344 155 346 157
rect 563 155 565 157
rect 611 155 613 157
rect 830 155 832 157
rect 37 143 39 145
rect 77 143 79 145
rect 296 143 298 145
rect 344 143 346 145
rect 563 143 565 145
rect 611 143 613 145
rect 830 143 832 145
rect 37 11 39 13
rect 77 11 79 13
rect 296 11 298 13
rect 344 11 346 13
rect 563 11 565 13
rect 611 11 613 13
rect 830 11 832 13
rect 460 -1 462 1
rect 698 -1 700 1
rect 460 -133 462 -131
rect 698 -133 700 -131
rect 460 -145 462 -143
rect 698 -145 700 -143
rect 460 -277 462 -275
rect 698 -277 700 -275
<< ptiect1 >>
rect 37 227 39 229
rect 77 227 79 229
rect 296 227 298 229
rect 344 227 346 229
rect 563 227 565 229
rect 611 227 613 229
rect 830 227 832 229
rect 37 215 39 217
rect 77 215 79 217
rect 296 215 298 217
rect 344 215 346 217
rect 563 215 565 217
rect 611 215 613 217
rect 830 215 832 217
rect 37 83 39 85
rect 77 83 79 85
rect 296 83 298 85
rect 344 83 346 85
rect 563 83 565 85
rect 611 83 613 85
rect 830 83 832 85
rect 37 71 39 73
rect 77 71 79 73
rect 296 71 298 73
rect 344 71 346 73
rect 563 71 565 73
rect 611 71 613 73
rect 830 71 832 73
rect 427 -61 429 -59
rect 698 -61 700 -59
rect 427 -73 429 -71
rect 698 -73 700 -71
rect 427 -205 429 -203
rect 698 -205 700 -203
rect 427 -217 429 -215
rect 698 -217 700 -215
<< pdifct0 >>
rect 8 277 10 279
rect 18 277 20 279
rect 18 270 20 272
rect 28 275 30 277
rect 48 277 50 279
rect 58 277 60 279
rect 58 270 60 272
rect 68 275 70 277
rect 99 284 101 286
rect 111 265 113 267
rect 134 284 136 286
rect 134 277 136 279
rect 146 276 148 278
rect 146 269 148 271
rect 156 284 158 286
rect 156 277 158 279
rect 188 284 190 286
rect 188 277 190 279
rect 198 276 200 278
rect 198 269 200 271
rect 210 284 212 286
rect 210 277 212 279
rect 245 284 247 286
rect 233 265 235 267
rect 267 277 269 279
rect 286 284 288 286
rect 315 277 317 279
rect 325 277 327 279
rect 325 270 327 272
rect 335 275 337 277
rect 366 284 368 286
rect 378 265 380 267
rect 401 284 403 286
rect 401 277 403 279
rect 413 276 415 278
rect 413 269 415 271
rect 423 284 425 286
rect 423 277 425 279
rect 455 284 457 286
rect 455 277 457 279
rect 465 276 467 278
rect 465 269 467 271
rect 477 284 479 286
rect 477 277 479 279
rect 512 284 514 286
rect 500 265 502 267
rect 534 277 536 279
rect 553 284 555 286
rect 582 277 584 279
rect 592 277 594 279
rect 592 270 594 272
rect 602 275 604 277
rect 633 284 635 286
rect 645 265 647 267
rect 668 284 670 286
rect 668 277 670 279
rect 680 276 682 278
rect 680 269 682 271
rect 690 284 692 286
rect 690 277 692 279
rect 722 284 724 286
rect 722 277 724 279
rect 732 276 734 278
rect 732 269 734 271
rect 744 284 746 286
rect 744 277 746 279
rect 779 284 781 286
rect 767 265 769 267
rect 801 277 803 279
rect 820 284 822 286
rect 8 165 10 167
rect 18 172 20 174
rect 18 165 20 167
rect 28 167 30 169
rect 48 165 50 167
rect 58 172 60 174
rect 58 165 60 167
rect 68 167 70 169
rect 111 177 113 179
rect 99 158 101 160
rect 134 165 136 167
rect 134 158 136 160
rect 146 173 148 175
rect 146 166 148 168
rect 156 165 158 167
rect 156 158 158 160
rect 188 165 190 167
rect 188 158 190 160
rect 198 173 200 175
rect 198 166 200 168
rect 210 165 212 167
rect 210 158 212 160
rect 233 177 235 179
rect 245 158 247 160
rect 267 165 269 167
rect 315 165 317 167
rect 325 172 327 174
rect 325 165 327 167
rect 335 167 337 169
rect 286 158 288 160
rect 378 177 380 179
rect 366 158 368 160
rect 401 165 403 167
rect 401 158 403 160
rect 413 173 415 175
rect 413 166 415 168
rect 423 165 425 167
rect 423 158 425 160
rect 455 165 457 167
rect 455 158 457 160
rect 465 173 467 175
rect 465 166 467 168
rect 477 165 479 167
rect 477 158 479 160
rect 500 177 502 179
rect 512 158 514 160
rect 534 165 536 167
rect 582 165 584 167
rect 592 172 594 174
rect 592 165 594 167
rect 602 167 604 169
rect 553 158 555 160
rect 645 177 647 179
rect 633 158 635 160
rect 668 165 670 167
rect 668 158 670 160
rect 680 173 682 175
rect 680 166 682 168
rect 690 165 692 167
rect 690 158 692 160
rect 722 165 724 167
rect 722 158 724 160
rect 732 173 734 175
rect 732 166 734 168
rect 744 165 746 167
rect 744 158 746 160
rect 767 177 769 179
rect 779 158 781 160
rect 801 165 803 167
rect 820 158 822 160
rect 8 133 10 135
rect 18 133 20 135
rect 18 126 20 128
rect 28 131 30 133
rect 48 133 50 135
rect 58 133 60 135
rect 58 126 60 128
rect 68 131 70 133
rect 99 140 101 142
rect 111 121 113 123
rect 134 140 136 142
rect 134 133 136 135
rect 146 132 148 134
rect 146 125 148 127
rect 156 140 158 142
rect 156 133 158 135
rect 188 140 190 142
rect 188 133 190 135
rect 198 132 200 134
rect 198 125 200 127
rect 210 140 212 142
rect 210 133 212 135
rect 245 140 247 142
rect 233 121 235 123
rect 267 133 269 135
rect 286 140 288 142
rect 315 133 317 135
rect 325 133 327 135
rect 325 126 327 128
rect 335 131 337 133
rect 366 140 368 142
rect 378 121 380 123
rect 401 140 403 142
rect 401 133 403 135
rect 413 132 415 134
rect 413 125 415 127
rect 423 140 425 142
rect 423 133 425 135
rect 455 140 457 142
rect 455 133 457 135
rect 465 132 467 134
rect 465 125 467 127
rect 477 140 479 142
rect 477 133 479 135
rect 512 140 514 142
rect 500 121 502 123
rect 534 133 536 135
rect 553 140 555 142
rect 582 133 584 135
rect 592 133 594 135
rect 592 126 594 128
rect 602 131 604 133
rect 633 140 635 142
rect 645 121 647 123
rect 668 140 670 142
rect 668 133 670 135
rect 680 132 682 134
rect 680 125 682 127
rect 690 140 692 142
rect 690 133 692 135
rect 722 140 724 142
rect 722 133 724 135
rect 732 132 734 134
rect 732 125 734 127
rect 744 140 746 142
rect 744 133 746 135
rect 779 140 781 142
rect 767 121 769 123
rect 801 133 803 135
rect 820 140 822 142
rect 8 21 10 23
rect 18 28 20 30
rect 18 21 20 23
rect 28 23 30 25
rect 48 21 50 23
rect 58 28 60 30
rect 58 21 60 23
rect 68 23 70 25
rect 111 33 113 35
rect 99 14 101 16
rect 134 21 136 23
rect 134 14 136 16
rect 146 29 148 31
rect 146 22 148 24
rect 156 21 158 23
rect 156 14 158 16
rect 188 21 190 23
rect 188 14 190 16
rect 198 29 200 31
rect 198 22 200 24
rect 210 21 212 23
rect 210 14 212 16
rect 233 33 235 35
rect 245 14 247 16
rect 267 21 269 23
rect 315 21 317 23
rect 325 28 327 30
rect 325 21 327 23
rect 335 23 337 25
rect 286 14 288 16
rect 378 33 380 35
rect 366 14 368 16
rect 401 21 403 23
rect 401 14 403 16
rect 413 29 415 31
rect 413 22 415 24
rect 423 21 425 23
rect 423 14 425 16
rect 455 21 457 23
rect 455 14 457 16
rect 465 29 467 31
rect 465 22 467 24
rect 477 21 479 23
rect 477 14 479 16
rect 500 33 502 35
rect 512 14 514 16
rect 534 21 536 23
rect 582 21 584 23
rect 592 28 594 30
rect 592 21 594 23
rect 602 23 604 25
rect 553 14 555 16
rect 645 33 647 35
rect 633 14 635 16
rect 668 21 670 23
rect 668 14 670 16
rect 680 29 682 31
rect 680 22 682 24
rect 690 21 692 23
rect 690 14 692 16
rect 722 21 724 23
rect 722 14 724 16
rect 732 29 734 31
rect 732 22 734 24
rect 744 21 746 23
rect 744 14 746 16
rect 767 33 769 35
rect 779 14 781 16
rect 801 21 803 23
rect 820 14 822 16
rect 434 -25 436 -23
rect 444 -4 446 -2
rect 444 -11 446 -9
rect 460 -18 462 -16
rect 460 -25 462 -23
rect 480 -10 482 -8
rect 501 -4 503 -2
rect 513 -23 515 -21
rect 536 -4 538 -2
rect 536 -11 538 -9
rect 548 -12 550 -10
rect 548 -19 550 -17
rect 558 -4 560 -2
rect 558 -11 560 -9
rect 590 -4 592 -2
rect 590 -11 592 -9
rect 600 -12 602 -10
rect 600 -19 602 -17
rect 612 -4 614 -2
rect 612 -11 614 -9
rect 647 -4 649 -2
rect 635 -23 637 -21
rect 669 -11 671 -9
rect 688 -4 690 -2
rect 722 -4 724 -2
rect 739 -14 741 -12
rect 756 -4 758 -2
rect 712 -26 714 -24
rect 786 -4 788 -2
rect 803 -14 805 -12
rect 820 -4 822 -2
rect 776 -26 778 -24
rect 434 -109 436 -107
rect 444 -123 446 -121
rect 460 -109 462 -107
rect 460 -116 462 -114
rect 444 -130 446 -128
rect 480 -124 482 -122
rect 513 -111 515 -109
rect 501 -130 503 -128
rect 536 -123 538 -121
rect 536 -130 538 -128
rect 548 -115 550 -113
rect 548 -122 550 -120
rect 558 -123 560 -121
rect 558 -130 560 -128
rect 590 -123 592 -121
rect 590 -130 592 -128
rect 600 -115 602 -113
rect 600 -122 602 -120
rect 612 -123 614 -121
rect 612 -130 614 -128
rect 635 -111 637 -109
rect 647 -130 649 -128
rect 669 -123 671 -121
rect 712 -108 714 -106
rect 776 -108 778 -106
rect 688 -130 690 -128
rect 722 -130 724 -128
rect 739 -120 741 -118
rect 756 -130 758 -128
rect 786 -130 788 -128
rect 803 -120 805 -118
rect 820 -130 822 -128
rect 434 -169 436 -167
rect 444 -148 446 -146
rect 444 -155 446 -153
rect 460 -162 462 -160
rect 460 -169 462 -167
rect 480 -154 482 -152
rect 501 -148 503 -146
rect 513 -167 515 -165
rect 536 -148 538 -146
rect 536 -155 538 -153
rect 548 -156 550 -154
rect 548 -163 550 -161
rect 558 -148 560 -146
rect 558 -155 560 -153
rect 590 -148 592 -146
rect 590 -155 592 -153
rect 600 -156 602 -154
rect 600 -163 602 -161
rect 612 -148 614 -146
rect 612 -155 614 -153
rect 647 -148 649 -146
rect 635 -167 637 -165
rect 669 -155 671 -153
rect 688 -148 690 -146
rect 722 -148 724 -146
rect 739 -158 741 -156
rect 756 -148 758 -146
rect 712 -170 714 -168
rect 786 -148 788 -146
rect 803 -158 805 -156
rect 820 -148 822 -146
rect 776 -170 778 -168
rect 434 -253 436 -251
rect 444 -267 446 -265
rect 460 -253 462 -251
rect 460 -260 462 -258
rect 444 -274 446 -272
rect 480 -268 482 -266
rect 513 -255 515 -253
rect 501 -274 503 -272
rect 536 -267 538 -265
rect 536 -274 538 -272
rect 548 -259 550 -257
rect 548 -266 550 -264
rect 558 -267 560 -265
rect 558 -274 560 -272
rect 590 -267 592 -265
rect 590 -274 592 -272
rect 600 -259 602 -257
rect 600 -266 602 -264
rect 612 -267 614 -265
rect 612 -274 614 -272
rect 635 -255 637 -253
rect 647 -274 649 -272
rect 669 -267 671 -265
rect 712 -252 714 -250
rect 776 -252 778 -250
rect 688 -274 690 -272
rect 722 -274 724 -272
rect 739 -264 741 -262
rect 756 -274 758 -272
rect 786 -274 788 -272
rect 803 -264 805 -262
rect 820 -274 822 -272
<< pdifct1 >>
rect 38 270 40 272
rect 38 263 40 265
rect 78 270 80 272
rect 78 263 80 265
rect 88 272 90 274
rect 88 265 90 267
rect 166 269 168 271
rect 166 262 168 264
rect 178 269 180 271
rect 178 262 180 264
rect 256 272 258 274
rect 256 265 258 267
rect 297 274 299 276
rect 297 267 299 269
rect 345 270 347 272
rect 345 263 347 265
rect 355 272 357 274
rect 355 265 357 267
rect 433 269 435 271
rect 433 262 435 264
rect 445 269 447 271
rect 445 262 447 264
rect 523 272 525 274
rect 523 265 525 267
rect 564 274 566 276
rect 564 267 566 269
rect 612 270 614 272
rect 612 263 614 265
rect 622 272 624 274
rect 622 265 624 267
rect 700 269 702 271
rect 700 262 702 264
rect 712 269 714 271
rect 712 262 714 264
rect 790 272 792 274
rect 790 265 792 267
rect 831 274 833 276
rect 831 267 833 269
rect 38 178 40 180
rect 38 170 40 172
rect 78 179 80 181
rect 78 172 80 174
rect 88 177 90 179
rect 88 170 90 172
rect 166 180 168 182
rect 166 173 168 175
rect 178 180 180 182
rect 178 173 180 175
rect 256 177 258 179
rect 256 170 258 172
rect 297 175 299 177
rect 297 168 299 170
rect 345 179 347 181
rect 345 172 347 174
rect 355 177 357 179
rect 355 170 357 172
rect 433 180 435 182
rect 433 173 435 175
rect 445 180 447 182
rect 445 173 447 175
rect 523 177 525 179
rect 523 170 525 172
rect 564 175 566 177
rect 564 168 566 170
rect 612 179 614 181
rect 612 172 614 174
rect 622 177 624 179
rect 622 170 624 172
rect 700 180 702 182
rect 700 173 702 175
rect 712 180 714 182
rect 712 173 714 175
rect 790 177 792 179
rect 790 170 792 172
rect 831 175 833 177
rect 831 168 833 170
rect 38 129 40 131
rect 38 121 40 123
rect 78 126 80 128
rect 78 119 80 121
rect 88 128 90 130
rect 88 121 90 123
rect 166 125 168 127
rect 166 118 168 120
rect 178 125 180 127
rect 178 118 180 120
rect 256 128 258 130
rect 256 121 258 123
rect 297 130 299 132
rect 297 123 299 125
rect 345 126 347 128
rect 345 119 347 121
rect 355 128 357 130
rect 355 121 357 123
rect 433 125 435 127
rect 433 118 435 120
rect 445 125 447 127
rect 445 118 447 120
rect 523 128 525 130
rect 523 121 525 123
rect 564 130 566 132
rect 564 123 566 125
rect 612 126 614 128
rect 612 119 614 121
rect 622 128 624 130
rect 622 121 624 123
rect 700 125 702 127
rect 700 118 702 120
rect 712 125 714 127
rect 712 118 714 120
rect 790 128 792 130
rect 790 121 792 123
rect 831 130 833 132
rect 831 123 833 125
rect 38 35 40 37
rect 38 28 40 30
rect 78 35 80 37
rect 78 28 80 30
rect 88 33 90 35
rect 88 26 90 28
rect 166 36 168 38
rect 166 29 168 31
rect 178 36 180 38
rect 178 29 180 31
rect 256 33 258 35
rect 256 26 258 28
rect 297 31 299 33
rect 297 24 299 26
rect 345 35 347 37
rect 345 28 347 30
rect 355 33 357 35
rect 355 26 357 28
rect 433 36 435 38
rect 433 29 435 31
rect 445 36 447 38
rect 445 29 447 31
rect 523 33 525 35
rect 523 26 525 28
rect 564 31 566 33
rect 564 24 566 26
rect 612 35 614 37
rect 612 28 614 30
rect 622 33 624 35
rect 622 26 624 28
rect 700 36 702 38
rect 700 29 702 31
rect 712 36 714 38
rect 712 29 714 31
rect 790 33 792 35
rect 790 26 792 28
rect 831 31 833 33
rect 831 24 833 26
rect 470 -18 472 -16
rect 490 -16 492 -14
rect 490 -23 492 -21
rect 568 -19 570 -17
rect 568 -26 570 -24
rect 580 -19 582 -17
rect 580 -26 582 -24
rect 658 -16 660 -14
rect 658 -23 660 -21
rect 699 -14 701 -12
rect 699 -21 701 -19
rect 766 -11 768 -9
rect 830 -11 832 -9
rect 470 -116 472 -114
rect 490 -111 492 -109
rect 490 -118 492 -116
rect 568 -108 570 -106
rect 568 -115 570 -113
rect 580 -108 582 -106
rect 580 -115 582 -113
rect 658 -111 660 -109
rect 658 -118 660 -116
rect 699 -113 701 -111
rect 699 -120 701 -118
rect 766 -123 768 -121
rect 830 -123 832 -121
rect 470 -162 472 -160
rect 490 -160 492 -158
rect 490 -167 492 -165
rect 568 -163 570 -161
rect 568 -170 570 -168
rect 580 -163 582 -161
rect 580 -170 582 -168
rect 658 -160 660 -158
rect 658 -167 660 -165
rect 699 -158 701 -156
rect 699 -165 701 -163
rect 766 -155 768 -153
rect 830 -155 832 -153
rect 470 -260 472 -258
rect 490 -255 492 -253
rect 490 -262 492 -260
rect 568 -252 570 -250
rect 568 -259 570 -257
rect 580 -252 582 -250
rect 580 -259 582 -257
rect 658 -255 660 -253
rect 658 -262 660 -260
rect 699 -257 701 -255
rect 699 -264 701 -262
rect 766 -267 768 -265
rect 830 -267 832 -265
<< alu0 >>
rect 6 279 12 286
rect 6 277 8 279
rect 10 277 12 279
rect 6 276 12 277
rect 17 279 21 281
rect 17 277 18 279
rect 20 277 21 279
rect 17 272 21 277
rect 26 277 32 286
rect 26 275 28 277
rect 30 275 32 277
rect 46 279 52 286
rect 46 277 48 279
rect 50 277 52 279
rect 46 276 52 277
rect 57 279 61 281
rect 57 277 58 279
rect 60 277 61 279
rect 26 274 32 275
rect 17 270 18 272
rect 20 271 21 272
rect 20 270 34 271
rect 17 267 34 270
rect 30 255 34 267
rect 30 253 31 255
rect 33 253 34 255
rect 30 248 34 253
rect 22 244 34 248
rect 57 272 61 277
rect 66 277 72 286
rect 97 284 99 286
rect 101 284 103 286
rect 97 283 103 284
rect 132 284 134 286
rect 136 284 138 286
rect 66 275 68 277
rect 70 275 72 277
rect 132 279 138 284
rect 154 284 156 286
rect 158 284 160 286
rect 132 277 134 279
rect 136 277 138 279
rect 132 276 138 277
rect 145 278 149 280
rect 145 276 146 278
rect 148 276 149 278
rect 154 279 160 284
rect 154 277 156 279
rect 158 277 160 279
rect 154 276 160 277
rect 186 284 188 286
rect 190 284 192 286
rect 186 279 192 284
rect 208 284 210 286
rect 212 284 214 286
rect 186 277 188 279
rect 190 277 192 279
rect 186 276 192 277
rect 197 278 201 280
rect 197 276 198 278
rect 200 276 201 278
rect 208 279 214 284
rect 243 284 245 286
rect 247 284 249 286
rect 243 283 249 284
rect 284 284 286 286
rect 288 284 290 286
rect 284 283 290 284
rect 208 277 210 279
rect 212 277 214 279
rect 208 276 214 277
rect 265 279 282 280
rect 265 277 267 279
rect 269 277 282 279
rect 265 276 282 277
rect 313 279 319 286
rect 313 277 315 279
rect 317 277 319 279
rect 313 276 319 277
rect 324 279 328 281
rect 324 277 325 279
rect 327 277 328 279
rect 66 274 72 275
rect 57 270 58 272
rect 60 271 61 272
rect 60 270 74 271
rect 57 267 74 270
rect 22 240 26 244
rect 37 241 38 243
rect 70 255 74 267
rect 70 253 71 255
rect 73 253 74 255
rect 70 248 74 253
rect 62 244 74 248
rect 6 239 26 240
rect 6 237 8 239
rect 10 237 26 239
rect 6 236 26 237
rect 62 240 66 244
rect 77 241 78 243
rect 46 239 66 240
rect 46 237 48 239
rect 50 237 66 239
rect 46 236 66 237
rect 102 272 126 276
rect 145 272 149 276
rect 100 268 106 272
rect 122 271 162 272
rect 122 269 146 271
rect 148 269 162 271
rect 100 258 104 268
rect 110 267 114 269
rect 122 268 162 269
rect 110 265 111 267
rect 113 265 114 267
rect 110 264 114 265
rect 100 256 101 258
rect 103 256 104 258
rect 100 254 104 256
rect 107 260 114 264
rect 107 249 111 260
rect 150 255 154 260
rect 150 253 151 255
rect 153 253 154 255
rect 93 248 111 249
rect 93 246 95 248
rect 97 247 111 248
rect 97 246 122 247
rect 93 245 118 246
rect 107 244 118 245
rect 120 244 122 246
rect 107 243 122 244
rect 127 246 131 248
rect 127 244 128 246
rect 130 244 131 246
rect 127 239 131 244
rect 150 251 154 253
rect 158 257 162 268
rect 158 255 164 257
rect 158 253 161 255
rect 163 253 164 255
rect 158 251 164 253
rect 158 248 162 251
rect 142 244 162 248
rect 142 240 146 244
rect 106 238 128 239
rect 97 235 101 237
rect 106 236 108 238
rect 110 237 128 238
rect 130 237 131 239
rect 110 236 131 237
rect 136 239 146 240
rect 136 237 138 239
rect 140 237 146 239
rect 136 236 146 237
rect 197 272 201 276
rect 220 272 244 276
rect 184 271 224 272
rect 184 269 198 271
rect 200 269 224 271
rect 184 268 224 269
rect 184 257 188 268
rect 232 267 236 269
rect 240 268 246 272
rect 232 265 233 267
rect 235 265 236 267
rect 232 264 236 265
rect 232 260 239 264
rect 182 255 188 257
rect 182 253 183 255
rect 185 253 188 255
rect 182 251 188 253
rect 192 255 196 260
rect 192 253 193 255
rect 195 253 196 255
rect 192 251 196 253
rect 184 248 188 251
rect 184 244 204 248
rect 200 240 204 244
rect 235 249 239 260
rect 242 258 246 268
rect 242 256 243 258
rect 245 256 246 258
rect 242 254 246 256
rect 235 248 253 249
rect 215 246 219 248
rect 235 247 249 248
rect 215 244 216 246
rect 218 244 219 246
rect 200 239 210 240
rect 200 237 206 239
rect 208 237 210 239
rect 200 236 210 237
rect 215 239 219 244
rect 224 246 249 247
rect 251 246 253 248
rect 224 244 226 246
rect 228 245 253 246
rect 228 244 239 245
rect 224 243 239 244
rect 278 272 282 276
rect 278 268 293 272
rect 268 259 274 260
rect 289 255 293 268
rect 296 265 297 276
rect 289 253 290 255
rect 292 253 293 255
rect 289 247 293 253
rect 324 272 328 277
rect 333 277 339 286
rect 364 284 366 286
rect 368 284 370 286
rect 364 283 370 284
rect 399 284 401 286
rect 403 284 405 286
rect 333 275 335 277
rect 337 275 339 277
rect 399 279 405 284
rect 421 284 423 286
rect 425 284 427 286
rect 399 277 401 279
rect 403 277 405 279
rect 399 276 405 277
rect 412 278 416 280
rect 412 276 413 278
rect 415 276 416 278
rect 421 279 427 284
rect 421 277 423 279
rect 425 277 427 279
rect 421 276 427 277
rect 453 284 455 286
rect 457 284 459 286
rect 453 279 459 284
rect 475 284 477 286
rect 479 284 481 286
rect 453 277 455 279
rect 457 277 459 279
rect 453 276 459 277
rect 464 278 468 280
rect 464 276 465 278
rect 467 276 468 278
rect 475 279 481 284
rect 510 284 512 286
rect 514 284 516 286
rect 510 283 516 284
rect 551 284 553 286
rect 555 284 557 286
rect 551 283 557 284
rect 475 277 477 279
rect 479 277 481 279
rect 475 276 481 277
rect 532 279 549 280
rect 532 277 534 279
rect 536 277 549 279
rect 532 276 549 277
rect 580 279 586 286
rect 580 277 582 279
rect 584 277 586 279
rect 580 276 586 277
rect 591 279 595 281
rect 591 277 592 279
rect 594 277 595 279
rect 333 274 339 275
rect 324 270 325 272
rect 327 271 328 272
rect 327 270 341 271
rect 324 267 341 270
rect 275 246 293 247
rect 275 244 277 246
rect 279 244 293 246
rect 275 243 293 244
rect 337 255 341 267
rect 337 253 338 255
rect 340 253 341 255
rect 337 248 341 253
rect 329 244 341 248
rect 329 240 333 244
rect 344 241 345 243
rect 215 237 216 239
rect 218 238 240 239
rect 218 237 236 238
rect 215 236 236 237
rect 238 236 240 238
rect 106 235 131 236
rect 215 235 240 236
rect 245 235 249 237
rect 313 239 333 240
rect 313 237 315 239
rect 317 237 333 239
rect 313 236 333 237
rect 369 272 393 276
rect 412 272 416 276
rect 367 268 373 272
rect 389 271 429 272
rect 389 269 413 271
rect 415 269 429 271
rect 367 258 371 268
rect 377 267 381 269
rect 389 268 429 269
rect 377 265 378 267
rect 380 265 381 267
rect 377 264 381 265
rect 367 256 368 258
rect 370 256 371 258
rect 367 254 371 256
rect 374 260 381 264
rect 374 249 378 260
rect 417 255 421 260
rect 417 253 418 255
rect 420 253 421 255
rect 360 248 378 249
rect 360 246 362 248
rect 364 247 378 248
rect 364 246 389 247
rect 360 245 385 246
rect 374 244 385 245
rect 387 244 389 246
rect 374 243 389 244
rect 394 246 398 248
rect 394 244 395 246
rect 397 244 398 246
rect 394 239 398 244
rect 417 251 421 253
rect 425 257 429 268
rect 425 255 431 257
rect 425 253 428 255
rect 430 253 431 255
rect 425 251 431 253
rect 425 248 429 251
rect 409 244 429 248
rect 409 240 413 244
rect 373 238 395 239
rect 364 235 368 237
rect 373 236 375 238
rect 377 237 395 238
rect 397 237 398 239
rect 377 236 398 237
rect 403 239 413 240
rect 403 237 405 239
rect 407 237 413 239
rect 403 236 413 237
rect 464 272 468 276
rect 487 272 511 276
rect 451 271 491 272
rect 451 269 465 271
rect 467 269 491 271
rect 451 268 491 269
rect 451 257 455 268
rect 499 267 503 269
rect 507 268 513 272
rect 499 265 500 267
rect 502 265 503 267
rect 499 264 503 265
rect 499 260 506 264
rect 449 255 455 257
rect 449 253 450 255
rect 452 253 455 255
rect 449 251 455 253
rect 459 255 463 260
rect 459 253 460 255
rect 462 253 463 255
rect 459 251 463 253
rect 451 248 455 251
rect 451 244 471 248
rect 467 240 471 244
rect 502 249 506 260
rect 509 258 513 268
rect 509 256 510 258
rect 512 256 513 258
rect 509 254 513 256
rect 502 248 520 249
rect 482 246 486 248
rect 502 247 516 248
rect 482 244 483 246
rect 485 244 486 246
rect 467 239 477 240
rect 467 237 473 239
rect 475 237 477 239
rect 467 236 477 237
rect 482 239 486 244
rect 491 246 516 247
rect 518 246 520 248
rect 491 244 493 246
rect 495 245 520 246
rect 545 272 549 276
rect 545 268 560 272
rect 535 259 541 260
rect 495 244 506 245
rect 491 243 506 244
rect 556 255 560 268
rect 563 265 564 276
rect 556 253 557 255
rect 559 253 560 255
rect 556 247 560 253
rect 591 272 595 277
rect 600 277 606 286
rect 631 284 633 286
rect 635 284 637 286
rect 631 283 637 284
rect 666 284 668 286
rect 670 284 672 286
rect 600 275 602 277
rect 604 275 606 277
rect 666 279 672 284
rect 688 284 690 286
rect 692 284 694 286
rect 666 277 668 279
rect 670 277 672 279
rect 666 276 672 277
rect 679 278 683 280
rect 679 276 680 278
rect 682 276 683 278
rect 688 279 694 284
rect 688 277 690 279
rect 692 277 694 279
rect 688 276 694 277
rect 720 284 722 286
rect 724 284 726 286
rect 720 279 726 284
rect 742 284 744 286
rect 746 284 748 286
rect 720 277 722 279
rect 724 277 726 279
rect 720 276 726 277
rect 731 278 735 280
rect 731 276 732 278
rect 734 276 735 278
rect 742 279 748 284
rect 777 284 779 286
rect 781 284 783 286
rect 777 283 783 284
rect 818 284 820 286
rect 822 284 824 286
rect 818 283 824 284
rect 742 277 744 279
rect 746 277 748 279
rect 742 276 748 277
rect 799 279 816 280
rect 799 277 801 279
rect 803 277 816 279
rect 799 276 816 277
rect 600 274 606 275
rect 591 270 592 272
rect 594 271 595 272
rect 594 270 608 271
rect 591 267 608 270
rect 542 246 560 247
rect 542 244 544 246
rect 546 244 560 246
rect 542 243 560 244
rect 604 255 608 267
rect 604 253 605 255
rect 607 253 608 255
rect 604 248 608 253
rect 596 244 608 248
rect 596 240 600 244
rect 611 241 612 243
rect 482 237 483 239
rect 485 238 507 239
rect 485 237 503 238
rect 482 236 503 237
rect 505 236 507 238
rect 373 235 398 236
rect 482 235 507 236
rect 512 235 516 237
rect 580 239 600 240
rect 580 237 582 239
rect 584 237 600 239
rect 580 236 600 237
rect 636 272 660 276
rect 679 272 683 276
rect 634 268 640 272
rect 656 271 696 272
rect 656 269 680 271
rect 682 269 696 271
rect 634 258 638 268
rect 644 267 648 269
rect 656 268 696 269
rect 644 265 645 267
rect 647 265 648 267
rect 644 264 648 265
rect 634 256 635 258
rect 637 256 638 258
rect 634 254 638 256
rect 641 260 648 264
rect 641 249 645 260
rect 684 255 688 260
rect 684 253 685 255
rect 687 253 688 255
rect 627 248 645 249
rect 627 246 629 248
rect 631 247 645 248
rect 631 246 656 247
rect 627 245 652 246
rect 641 244 652 245
rect 654 244 656 246
rect 641 243 656 244
rect 661 246 665 248
rect 661 244 662 246
rect 664 244 665 246
rect 661 239 665 244
rect 684 251 688 253
rect 692 257 696 268
rect 692 255 698 257
rect 692 253 695 255
rect 697 253 698 255
rect 692 251 698 253
rect 692 248 696 251
rect 676 244 696 248
rect 676 240 680 244
rect 640 238 662 239
rect 631 235 635 237
rect 640 236 642 238
rect 644 237 662 238
rect 664 237 665 239
rect 644 236 665 237
rect 670 239 680 240
rect 670 237 672 239
rect 674 237 680 239
rect 670 236 680 237
rect 731 272 735 276
rect 754 272 778 276
rect 718 271 758 272
rect 718 269 732 271
rect 734 269 758 271
rect 718 268 758 269
rect 718 257 722 268
rect 766 267 770 269
rect 774 268 780 272
rect 766 265 767 267
rect 769 265 770 267
rect 766 264 770 265
rect 766 260 773 264
rect 716 255 722 257
rect 716 253 717 255
rect 719 253 722 255
rect 716 251 722 253
rect 726 255 730 260
rect 726 253 727 255
rect 729 253 730 255
rect 726 251 730 253
rect 718 248 722 251
rect 718 244 738 248
rect 734 240 738 244
rect 769 249 773 260
rect 776 258 780 268
rect 776 256 777 258
rect 779 256 780 258
rect 776 254 780 256
rect 769 248 787 249
rect 749 246 753 248
rect 769 247 783 248
rect 749 244 750 246
rect 752 244 753 246
rect 734 239 744 240
rect 734 237 740 239
rect 742 237 744 239
rect 734 236 744 237
rect 749 239 753 244
rect 758 246 783 247
rect 785 246 787 248
rect 758 244 760 246
rect 762 245 787 246
rect 812 272 816 276
rect 812 268 827 272
rect 802 259 808 260
rect 762 244 773 245
rect 758 243 773 244
rect 823 255 827 268
rect 830 265 831 276
rect 823 253 824 255
rect 826 253 827 255
rect 823 247 827 253
rect 809 246 827 247
rect 809 244 811 246
rect 813 244 827 246
rect 809 243 827 244
rect 749 237 750 239
rect 752 238 774 239
rect 752 237 770 238
rect 749 236 770 237
rect 772 236 774 238
rect 640 235 665 236
rect 749 235 774 236
rect 779 235 783 237
rect 97 233 98 235
rect 100 233 101 235
rect 245 233 246 235
rect 248 233 249 235
rect 97 230 101 233
rect 153 232 159 233
rect 153 230 155 232
rect 157 230 159 232
rect 187 232 193 233
rect 187 230 189 232
rect 191 230 193 232
rect 245 230 249 233
rect 265 233 271 234
rect 265 231 267 233
rect 269 231 271 233
rect 265 230 271 231
rect 284 233 290 234
rect 284 231 286 233
rect 288 231 290 233
rect 284 230 290 231
rect 364 233 365 235
rect 367 233 368 235
rect 512 233 513 235
rect 515 233 516 235
rect 364 230 368 233
rect 420 232 426 233
rect 420 230 422 232
rect 424 230 426 232
rect 454 232 460 233
rect 454 230 456 232
rect 458 230 460 232
rect 512 230 516 233
rect 532 233 538 234
rect 532 231 534 233
rect 536 231 538 233
rect 532 230 538 231
rect 551 233 557 234
rect 551 231 553 233
rect 555 231 557 233
rect 551 230 557 231
rect 631 233 632 235
rect 634 233 635 235
rect 779 233 780 235
rect 782 233 783 235
rect 631 230 635 233
rect 687 232 693 233
rect 687 230 689 232
rect 691 230 693 232
rect 721 232 727 233
rect 721 230 723 232
rect 725 230 727 232
rect 779 230 783 233
rect 799 233 805 234
rect 799 231 801 233
rect 803 231 805 233
rect 799 230 805 231
rect 818 233 824 234
rect 818 231 820 233
rect 822 231 824 233
rect 818 230 824 231
rect 97 211 101 214
rect 153 212 155 214
rect 157 212 159 214
rect 153 211 159 212
rect 187 212 189 214
rect 191 212 193 214
rect 187 211 193 212
rect 245 211 249 214
rect 97 209 98 211
rect 100 209 101 211
rect 245 209 246 211
rect 248 209 249 211
rect 265 213 271 214
rect 265 211 267 213
rect 269 211 271 213
rect 265 210 271 211
rect 284 213 290 214
rect 284 211 286 213
rect 288 211 290 213
rect 284 210 290 211
rect 364 211 368 214
rect 420 212 422 214
rect 424 212 426 214
rect 420 211 426 212
rect 454 212 456 214
rect 458 212 460 214
rect 454 211 460 212
rect 512 211 516 214
rect 364 209 365 211
rect 367 209 368 211
rect 512 209 513 211
rect 515 209 516 211
rect 532 213 538 214
rect 532 211 534 213
rect 536 211 538 213
rect 532 210 538 211
rect 551 213 557 214
rect 551 211 553 213
rect 555 211 557 213
rect 551 210 557 211
rect 631 211 635 214
rect 687 212 689 214
rect 691 212 693 214
rect 687 211 693 212
rect 721 212 723 214
rect 725 212 727 214
rect 721 211 727 212
rect 779 211 783 214
rect 631 209 632 211
rect 634 209 635 211
rect 779 209 780 211
rect 782 209 783 211
rect 799 213 805 214
rect 799 211 801 213
rect 803 211 805 213
rect 799 210 805 211
rect 818 213 824 214
rect 818 211 820 213
rect 822 211 824 213
rect 818 210 824 211
rect 6 207 26 208
rect 6 205 8 207
rect 10 205 26 207
rect 6 204 26 205
rect 22 200 26 204
rect 46 207 66 208
rect 46 205 48 207
rect 50 205 66 207
rect 46 204 66 205
rect 37 201 38 203
rect 22 196 34 200
rect 30 191 34 196
rect 30 189 31 191
rect 33 189 34 191
rect 30 177 34 189
rect 62 200 66 204
rect 77 201 78 203
rect 62 196 74 200
rect 70 191 74 196
rect 70 189 71 191
rect 73 189 74 191
rect 17 174 34 177
rect 17 172 18 174
rect 20 173 34 174
rect 20 172 21 173
rect 6 167 12 168
rect 6 165 8 167
rect 10 165 12 167
rect 6 158 12 165
rect 17 167 21 172
rect 70 177 74 189
rect 57 174 74 177
rect 57 172 58 174
rect 60 173 74 174
rect 60 172 61 173
rect 17 165 18 167
rect 20 165 21 167
rect 17 163 21 165
rect 26 169 32 170
rect 26 167 28 169
rect 30 167 32 169
rect 26 158 32 167
rect 46 167 52 168
rect 46 165 48 167
rect 50 165 52 167
rect 46 158 52 165
rect 57 167 61 172
rect 97 207 101 209
rect 106 208 131 209
rect 215 208 240 209
rect 106 206 108 208
rect 110 207 131 208
rect 110 206 128 207
rect 106 205 128 206
rect 130 205 131 207
rect 107 200 122 201
rect 107 199 118 200
rect 93 198 118 199
rect 120 198 122 200
rect 93 196 95 198
rect 97 197 122 198
rect 127 200 131 205
rect 136 207 146 208
rect 136 205 138 207
rect 140 205 146 207
rect 136 204 146 205
rect 127 198 128 200
rect 130 198 131 200
rect 97 196 111 197
rect 127 196 131 198
rect 93 195 111 196
rect 100 188 104 190
rect 100 186 101 188
rect 103 186 104 188
rect 100 176 104 186
rect 107 184 111 195
rect 142 200 146 204
rect 142 196 162 200
rect 158 193 162 196
rect 150 191 154 193
rect 150 189 151 191
rect 153 189 154 191
rect 150 184 154 189
rect 158 191 164 193
rect 158 189 161 191
rect 163 189 164 191
rect 158 187 164 189
rect 107 180 114 184
rect 110 179 114 180
rect 110 177 111 179
rect 113 177 114 179
rect 100 172 106 176
rect 110 175 114 177
rect 158 176 162 187
rect 122 175 162 176
rect 122 173 146 175
rect 148 173 162 175
rect 122 172 162 173
rect 57 165 58 167
rect 60 165 61 167
rect 57 163 61 165
rect 66 169 72 170
rect 66 167 68 169
rect 70 167 72 169
rect 102 168 126 172
rect 145 168 149 172
rect 200 207 210 208
rect 200 205 206 207
rect 208 205 210 207
rect 200 204 210 205
rect 215 207 236 208
rect 215 205 216 207
rect 218 206 236 207
rect 238 206 240 208
rect 245 207 249 209
rect 218 205 240 206
rect 200 200 204 204
rect 184 196 204 200
rect 184 193 188 196
rect 182 191 188 193
rect 182 189 183 191
rect 185 189 188 191
rect 182 187 188 189
rect 184 176 188 187
rect 192 191 196 193
rect 215 200 219 205
rect 313 207 333 208
rect 313 205 315 207
rect 317 205 333 207
rect 313 204 333 205
rect 215 198 216 200
rect 218 198 219 200
rect 215 196 219 198
rect 224 200 239 201
rect 224 198 226 200
rect 228 199 239 200
rect 228 198 253 199
rect 224 197 249 198
rect 235 196 249 197
rect 251 196 253 198
rect 235 195 253 196
rect 192 189 193 191
rect 195 189 196 191
rect 192 184 196 189
rect 235 184 239 195
rect 232 180 239 184
rect 242 188 246 190
rect 242 186 243 188
rect 245 186 246 188
rect 232 179 236 180
rect 232 177 233 179
rect 235 177 236 179
rect 184 175 224 176
rect 232 175 236 177
rect 242 176 246 186
rect 275 200 293 201
rect 275 198 277 200
rect 279 198 293 200
rect 275 197 293 198
rect 289 191 293 197
rect 289 189 290 191
rect 292 189 293 191
rect 268 184 274 185
rect 184 173 198 175
rect 200 173 224 175
rect 184 172 224 173
rect 240 172 246 176
rect 197 168 201 172
rect 220 168 244 172
rect 289 176 293 189
rect 278 172 293 176
rect 278 168 282 172
rect 296 168 297 179
rect 329 200 333 204
rect 344 201 345 203
rect 329 196 341 200
rect 337 191 341 196
rect 337 189 338 191
rect 340 189 341 191
rect 337 177 341 189
rect 324 174 341 177
rect 324 172 325 174
rect 327 173 341 174
rect 327 172 328 173
rect 66 158 72 167
rect 132 167 138 168
rect 132 165 134 167
rect 136 165 138 167
rect 97 160 103 161
rect 97 158 99 160
rect 101 158 103 160
rect 132 160 138 165
rect 145 166 146 168
rect 148 166 149 168
rect 145 164 149 166
rect 154 167 160 168
rect 154 165 156 167
rect 158 165 160 167
rect 132 158 134 160
rect 136 158 138 160
rect 154 160 160 165
rect 154 158 156 160
rect 158 158 160 160
rect 186 167 192 168
rect 186 165 188 167
rect 190 165 192 167
rect 186 160 192 165
rect 197 166 198 168
rect 200 166 201 168
rect 197 164 201 166
rect 208 167 214 168
rect 208 165 210 167
rect 212 165 214 167
rect 186 158 188 160
rect 190 158 192 160
rect 208 160 214 165
rect 265 167 282 168
rect 265 165 267 167
rect 269 165 282 167
rect 265 164 282 165
rect 313 167 319 168
rect 313 165 315 167
rect 317 165 319 167
rect 208 158 210 160
rect 212 158 214 160
rect 243 160 249 161
rect 243 158 245 160
rect 247 158 249 160
rect 284 160 290 161
rect 284 158 286 160
rect 288 158 290 160
rect 313 158 319 165
rect 324 167 328 172
rect 364 207 368 209
rect 373 208 398 209
rect 482 208 507 209
rect 373 206 375 208
rect 377 207 398 208
rect 377 206 395 207
rect 373 205 395 206
rect 397 205 398 207
rect 374 200 389 201
rect 374 199 385 200
rect 360 198 385 199
rect 387 198 389 200
rect 360 196 362 198
rect 364 197 389 198
rect 394 200 398 205
rect 403 207 413 208
rect 403 205 405 207
rect 407 205 413 207
rect 403 204 413 205
rect 394 198 395 200
rect 397 198 398 200
rect 364 196 378 197
rect 394 196 398 198
rect 360 195 378 196
rect 367 188 371 190
rect 367 186 368 188
rect 370 186 371 188
rect 367 176 371 186
rect 374 184 378 195
rect 409 200 413 204
rect 409 196 429 200
rect 425 193 429 196
rect 417 191 421 193
rect 417 189 418 191
rect 420 189 421 191
rect 417 184 421 189
rect 425 191 431 193
rect 425 189 428 191
rect 430 189 431 191
rect 425 187 431 189
rect 374 180 381 184
rect 377 179 381 180
rect 377 177 378 179
rect 380 177 381 179
rect 367 172 373 176
rect 377 175 381 177
rect 425 176 429 187
rect 389 175 429 176
rect 389 173 413 175
rect 415 173 429 175
rect 389 172 429 173
rect 324 165 325 167
rect 327 165 328 167
rect 324 163 328 165
rect 333 169 339 170
rect 333 167 335 169
rect 337 167 339 169
rect 369 168 393 172
rect 412 168 416 172
rect 467 207 477 208
rect 467 205 473 207
rect 475 205 477 207
rect 467 204 477 205
rect 482 207 503 208
rect 482 205 483 207
rect 485 206 503 207
rect 505 206 507 208
rect 512 207 516 209
rect 485 205 507 206
rect 467 200 471 204
rect 451 196 471 200
rect 451 193 455 196
rect 449 191 455 193
rect 449 189 450 191
rect 452 189 455 191
rect 449 187 455 189
rect 451 176 455 187
rect 459 191 463 193
rect 482 200 486 205
rect 580 207 600 208
rect 580 205 582 207
rect 584 205 600 207
rect 580 204 600 205
rect 482 198 483 200
rect 485 198 486 200
rect 482 196 486 198
rect 491 200 506 201
rect 491 198 493 200
rect 495 199 506 200
rect 495 198 520 199
rect 491 197 516 198
rect 502 196 516 197
rect 518 196 520 198
rect 502 195 520 196
rect 459 189 460 191
rect 462 189 463 191
rect 459 184 463 189
rect 502 184 506 195
rect 499 180 506 184
rect 509 188 513 190
rect 509 186 510 188
rect 512 186 513 188
rect 499 179 503 180
rect 499 177 500 179
rect 502 177 503 179
rect 451 175 491 176
rect 499 175 503 177
rect 509 176 513 186
rect 542 200 560 201
rect 542 198 544 200
rect 546 198 560 200
rect 542 197 560 198
rect 556 191 560 197
rect 556 189 557 191
rect 559 189 560 191
rect 535 184 541 185
rect 451 173 465 175
rect 467 173 491 175
rect 451 172 491 173
rect 507 172 513 176
rect 464 168 468 172
rect 487 168 511 172
rect 556 176 560 189
rect 545 172 560 176
rect 545 168 549 172
rect 563 168 564 179
rect 596 200 600 204
rect 611 201 612 203
rect 596 196 608 200
rect 604 191 608 196
rect 604 189 605 191
rect 607 189 608 191
rect 604 177 608 189
rect 591 174 608 177
rect 591 172 592 174
rect 594 173 608 174
rect 594 172 595 173
rect 333 158 339 167
rect 399 167 405 168
rect 399 165 401 167
rect 403 165 405 167
rect 364 160 370 161
rect 364 158 366 160
rect 368 158 370 160
rect 399 160 405 165
rect 412 166 413 168
rect 415 166 416 168
rect 412 164 416 166
rect 421 167 427 168
rect 421 165 423 167
rect 425 165 427 167
rect 399 158 401 160
rect 403 158 405 160
rect 421 160 427 165
rect 421 158 423 160
rect 425 158 427 160
rect 453 167 459 168
rect 453 165 455 167
rect 457 165 459 167
rect 453 160 459 165
rect 464 166 465 168
rect 467 166 468 168
rect 464 164 468 166
rect 475 167 481 168
rect 475 165 477 167
rect 479 165 481 167
rect 453 158 455 160
rect 457 158 459 160
rect 475 160 481 165
rect 532 167 549 168
rect 532 165 534 167
rect 536 165 549 167
rect 532 164 549 165
rect 580 167 586 168
rect 580 165 582 167
rect 584 165 586 167
rect 475 158 477 160
rect 479 158 481 160
rect 510 160 516 161
rect 510 158 512 160
rect 514 158 516 160
rect 551 160 557 161
rect 551 158 553 160
rect 555 158 557 160
rect 580 158 586 165
rect 591 167 595 172
rect 631 207 635 209
rect 640 208 665 209
rect 749 208 774 209
rect 640 206 642 208
rect 644 207 665 208
rect 644 206 662 207
rect 640 205 662 206
rect 664 205 665 207
rect 641 200 656 201
rect 641 199 652 200
rect 627 198 652 199
rect 654 198 656 200
rect 627 196 629 198
rect 631 197 656 198
rect 661 200 665 205
rect 670 207 680 208
rect 670 205 672 207
rect 674 205 680 207
rect 670 204 680 205
rect 661 198 662 200
rect 664 198 665 200
rect 631 196 645 197
rect 661 196 665 198
rect 627 195 645 196
rect 634 188 638 190
rect 634 186 635 188
rect 637 186 638 188
rect 634 176 638 186
rect 641 184 645 195
rect 676 200 680 204
rect 676 196 696 200
rect 692 193 696 196
rect 684 191 688 193
rect 684 189 685 191
rect 687 189 688 191
rect 684 184 688 189
rect 692 191 698 193
rect 692 189 695 191
rect 697 189 698 191
rect 692 187 698 189
rect 641 180 648 184
rect 644 179 648 180
rect 644 177 645 179
rect 647 177 648 179
rect 634 172 640 176
rect 644 175 648 177
rect 692 176 696 187
rect 656 175 696 176
rect 656 173 680 175
rect 682 173 696 175
rect 656 172 696 173
rect 591 165 592 167
rect 594 165 595 167
rect 591 163 595 165
rect 600 169 606 170
rect 600 167 602 169
rect 604 167 606 169
rect 636 168 660 172
rect 679 168 683 172
rect 734 207 744 208
rect 734 205 740 207
rect 742 205 744 207
rect 734 204 744 205
rect 749 207 770 208
rect 749 205 750 207
rect 752 206 770 207
rect 772 206 774 208
rect 779 207 783 209
rect 752 205 774 206
rect 734 200 738 204
rect 718 196 738 200
rect 718 193 722 196
rect 716 191 722 193
rect 716 189 717 191
rect 719 189 722 191
rect 716 187 722 189
rect 718 176 722 187
rect 726 191 730 193
rect 749 200 753 205
rect 749 198 750 200
rect 752 198 753 200
rect 749 196 753 198
rect 758 200 773 201
rect 758 198 760 200
rect 762 199 773 200
rect 762 198 787 199
rect 758 197 783 198
rect 769 196 783 197
rect 785 196 787 198
rect 769 195 787 196
rect 726 189 727 191
rect 729 189 730 191
rect 726 184 730 189
rect 769 184 773 195
rect 766 180 773 184
rect 776 188 780 190
rect 776 186 777 188
rect 779 186 780 188
rect 766 179 770 180
rect 766 177 767 179
rect 769 177 770 179
rect 718 175 758 176
rect 766 175 770 177
rect 776 176 780 186
rect 809 200 827 201
rect 809 198 811 200
rect 813 198 827 200
rect 809 197 827 198
rect 823 191 827 197
rect 823 189 824 191
rect 826 189 827 191
rect 802 184 808 185
rect 718 173 732 175
rect 734 173 758 175
rect 718 172 758 173
rect 774 172 780 176
rect 731 168 735 172
rect 754 168 778 172
rect 823 176 827 189
rect 812 172 827 176
rect 812 168 816 172
rect 830 168 831 179
rect 600 158 606 167
rect 666 167 672 168
rect 666 165 668 167
rect 670 165 672 167
rect 631 160 637 161
rect 631 158 633 160
rect 635 158 637 160
rect 666 160 672 165
rect 679 166 680 168
rect 682 166 683 168
rect 679 164 683 166
rect 688 167 694 168
rect 688 165 690 167
rect 692 165 694 167
rect 666 158 668 160
rect 670 158 672 160
rect 688 160 694 165
rect 688 158 690 160
rect 692 158 694 160
rect 720 167 726 168
rect 720 165 722 167
rect 724 165 726 167
rect 720 160 726 165
rect 731 166 732 168
rect 734 166 735 168
rect 731 164 735 166
rect 742 167 748 168
rect 742 165 744 167
rect 746 165 748 167
rect 720 158 722 160
rect 724 158 726 160
rect 742 160 748 165
rect 799 167 816 168
rect 799 165 801 167
rect 803 165 816 167
rect 799 164 816 165
rect 742 158 744 160
rect 746 158 748 160
rect 777 160 783 161
rect 777 158 779 160
rect 781 158 783 160
rect 818 160 824 161
rect 818 158 820 160
rect 822 158 824 160
rect 6 135 12 142
rect 6 133 8 135
rect 10 133 12 135
rect 6 132 12 133
rect 17 135 21 137
rect 17 133 18 135
rect 20 133 21 135
rect 17 128 21 133
rect 26 133 32 142
rect 46 135 52 142
rect 46 133 48 135
rect 50 133 52 135
rect 26 131 28 133
rect 30 131 32 133
rect 26 130 32 131
rect 46 132 52 133
rect 57 135 61 137
rect 57 133 58 135
rect 60 133 61 135
rect 17 126 18 128
rect 20 127 21 128
rect 20 126 34 127
rect 17 123 34 126
rect 30 111 34 123
rect 57 128 61 133
rect 66 133 72 142
rect 97 140 99 142
rect 101 140 103 142
rect 97 139 103 140
rect 132 140 134 142
rect 136 140 138 142
rect 66 131 68 133
rect 70 131 72 133
rect 132 135 138 140
rect 154 140 156 142
rect 158 140 160 142
rect 132 133 134 135
rect 136 133 138 135
rect 132 132 138 133
rect 145 134 149 136
rect 145 132 146 134
rect 148 132 149 134
rect 154 135 160 140
rect 154 133 156 135
rect 158 133 160 135
rect 154 132 160 133
rect 186 140 188 142
rect 190 140 192 142
rect 186 135 192 140
rect 208 140 210 142
rect 212 140 214 142
rect 186 133 188 135
rect 190 133 192 135
rect 186 132 192 133
rect 197 134 201 136
rect 197 132 198 134
rect 200 132 201 134
rect 208 135 214 140
rect 243 140 245 142
rect 247 140 249 142
rect 243 139 249 140
rect 284 140 286 142
rect 288 140 290 142
rect 284 139 290 140
rect 208 133 210 135
rect 212 133 214 135
rect 208 132 214 133
rect 265 135 282 136
rect 265 133 267 135
rect 269 133 282 135
rect 265 132 282 133
rect 313 135 319 142
rect 313 133 315 135
rect 317 133 319 135
rect 313 132 319 133
rect 324 135 328 137
rect 324 133 325 135
rect 327 133 328 135
rect 66 130 72 131
rect 57 126 58 128
rect 60 127 61 128
rect 60 126 74 127
rect 57 123 74 126
rect 30 109 31 111
rect 33 109 34 111
rect 30 104 34 109
rect 22 100 34 104
rect 22 96 26 100
rect 37 97 38 99
rect 70 111 74 123
rect 70 109 71 111
rect 73 109 74 111
rect 70 104 74 109
rect 62 100 74 104
rect 6 95 26 96
rect 6 93 8 95
rect 10 93 26 95
rect 6 92 26 93
rect 62 96 66 100
rect 77 97 78 99
rect 46 95 66 96
rect 46 93 48 95
rect 50 93 66 95
rect 46 92 66 93
rect 102 128 126 132
rect 145 128 149 132
rect 100 124 106 128
rect 122 127 162 128
rect 122 125 146 127
rect 148 125 162 127
rect 100 114 104 124
rect 110 123 114 125
rect 122 124 162 125
rect 110 121 111 123
rect 113 121 114 123
rect 110 120 114 121
rect 100 112 101 114
rect 103 112 104 114
rect 100 110 104 112
rect 107 116 114 120
rect 107 105 111 116
rect 150 111 154 116
rect 150 109 151 111
rect 153 109 154 111
rect 93 104 111 105
rect 93 102 95 104
rect 97 103 111 104
rect 97 102 122 103
rect 93 101 118 102
rect 107 100 118 101
rect 120 100 122 102
rect 107 99 122 100
rect 127 102 131 104
rect 127 100 128 102
rect 130 100 131 102
rect 127 95 131 100
rect 150 107 154 109
rect 158 113 162 124
rect 158 111 164 113
rect 158 109 161 111
rect 163 109 164 111
rect 158 107 164 109
rect 158 104 162 107
rect 142 100 162 104
rect 142 96 146 100
rect 106 94 128 95
rect 97 91 101 93
rect 106 92 108 94
rect 110 93 128 94
rect 130 93 131 95
rect 110 92 131 93
rect 136 95 146 96
rect 136 93 138 95
rect 140 93 146 95
rect 136 92 146 93
rect 197 128 201 132
rect 220 128 244 132
rect 184 127 224 128
rect 184 125 198 127
rect 200 125 224 127
rect 184 124 224 125
rect 184 113 188 124
rect 232 123 236 125
rect 240 124 246 128
rect 232 121 233 123
rect 235 121 236 123
rect 232 120 236 121
rect 232 116 239 120
rect 182 111 188 113
rect 182 109 183 111
rect 185 109 188 111
rect 182 107 188 109
rect 192 111 196 116
rect 192 109 193 111
rect 195 109 196 111
rect 192 107 196 109
rect 184 104 188 107
rect 184 100 204 104
rect 200 96 204 100
rect 235 105 239 116
rect 242 114 246 124
rect 242 112 243 114
rect 245 112 246 114
rect 242 110 246 112
rect 235 104 253 105
rect 215 102 219 104
rect 235 103 249 104
rect 215 100 216 102
rect 218 100 219 102
rect 200 95 210 96
rect 200 93 206 95
rect 208 93 210 95
rect 200 92 210 93
rect 215 95 219 100
rect 224 102 249 103
rect 251 102 253 104
rect 224 100 226 102
rect 228 101 253 102
rect 228 100 239 101
rect 224 99 239 100
rect 278 128 282 132
rect 278 124 293 128
rect 268 115 274 116
rect 289 111 293 124
rect 296 121 297 132
rect 289 109 290 111
rect 292 109 293 111
rect 289 103 293 109
rect 324 128 328 133
rect 333 133 339 142
rect 364 140 366 142
rect 368 140 370 142
rect 364 139 370 140
rect 399 140 401 142
rect 403 140 405 142
rect 333 131 335 133
rect 337 131 339 133
rect 399 135 405 140
rect 421 140 423 142
rect 425 140 427 142
rect 399 133 401 135
rect 403 133 405 135
rect 399 132 405 133
rect 412 134 416 136
rect 412 132 413 134
rect 415 132 416 134
rect 421 135 427 140
rect 421 133 423 135
rect 425 133 427 135
rect 421 132 427 133
rect 453 140 455 142
rect 457 140 459 142
rect 453 135 459 140
rect 475 140 477 142
rect 479 140 481 142
rect 453 133 455 135
rect 457 133 459 135
rect 453 132 459 133
rect 464 134 468 136
rect 464 132 465 134
rect 467 132 468 134
rect 475 135 481 140
rect 510 140 512 142
rect 514 140 516 142
rect 510 139 516 140
rect 551 140 553 142
rect 555 140 557 142
rect 551 139 557 140
rect 475 133 477 135
rect 479 133 481 135
rect 475 132 481 133
rect 532 135 549 136
rect 532 133 534 135
rect 536 133 549 135
rect 532 132 549 133
rect 580 135 586 142
rect 580 133 582 135
rect 584 133 586 135
rect 580 132 586 133
rect 591 135 595 137
rect 591 133 592 135
rect 594 133 595 135
rect 333 130 339 131
rect 324 126 325 128
rect 327 127 328 128
rect 327 126 341 127
rect 324 123 341 126
rect 275 102 293 103
rect 275 100 277 102
rect 279 100 293 102
rect 275 99 293 100
rect 337 111 341 123
rect 337 109 338 111
rect 340 109 341 111
rect 337 104 341 109
rect 329 100 341 104
rect 329 96 333 100
rect 344 97 345 99
rect 215 93 216 95
rect 218 94 240 95
rect 218 93 236 94
rect 215 92 236 93
rect 238 92 240 94
rect 106 91 131 92
rect 215 91 240 92
rect 245 91 249 93
rect 313 95 333 96
rect 313 93 315 95
rect 317 93 333 95
rect 313 92 333 93
rect 369 128 393 132
rect 412 128 416 132
rect 367 124 373 128
rect 389 127 429 128
rect 389 125 413 127
rect 415 125 429 127
rect 367 114 371 124
rect 377 123 381 125
rect 389 124 429 125
rect 377 121 378 123
rect 380 121 381 123
rect 377 120 381 121
rect 367 112 368 114
rect 370 112 371 114
rect 367 110 371 112
rect 374 116 381 120
rect 374 105 378 116
rect 417 111 421 116
rect 417 109 418 111
rect 420 109 421 111
rect 360 104 378 105
rect 360 102 362 104
rect 364 103 378 104
rect 364 102 389 103
rect 360 101 385 102
rect 374 100 385 101
rect 387 100 389 102
rect 374 99 389 100
rect 394 102 398 104
rect 394 100 395 102
rect 397 100 398 102
rect 394 95 398 100
rect 417 107 421 109
rect 425 113 429 124
rect 425 111 431 113
rect 425 109 428 111
rect 430 109 431 111
rect 425 107 431 109
rect 425 104 429 107
rect 409 100 429 104
rect 409 96 413 100
rect 373 94 395 95
rect 364 91 368 93
rect 373 92 375 94
rect 377 93 395 94
rect 397 93 398 95
rect 377 92 398 93
rect 403 95 413 96
rect 403 93 405 95
rect 407 93 413 95
rect 403 92 413 93
rect 464 128 468 132
rect 487 128 511 132
rect 451 127 491 128
rect 451 125 465 127
rect 467 125 491 127
rect 451 124 491 125
rect 451 113 455 124
rect 499 123 503 125
rect 507 124 513 128
rect 499 121 500 123
rect 502 121 503 123
rect 499 120 503 121
rect 499 116 506 120
rect 449 111 455 113
rect 449 109 450 111
rect 452 109 455 111
rect 449 107 455 109
rect 459 111 463 116
rect 459 109 460 111
rect 462 109 463 111
rect 459 107 463 109
rect 451 104 455 107
rect 451 100 471 104
rect 467 96 471 100
rect 502 105 506 116
rect 509 114 513 124
rect 509 112 510 114
rect 512 112 513 114
rect 509 110 513 112
rect 502 104 520 105
rect 482 102 486 104
rect 502 103 516 104
rect 482 100 483 102
rect 485 100 486 102
rect 467 95 477 96
rect 467 93 473 95
rect 475 93 477 95
rect 467 92 477 93
rect 482 95 486 100
rect 491 102 516 103
rect 518 102 520 104
rect 491 100 493 102
rect 495 101 520 102
rect 495 100 506 101
rect 491 99 506 100
rect 545 128 549 132
rect 545 124 560 128
rect 535 115 541 116
rect 556 111 560 124
rect 563 121 564 132
rect 556 109 557 111
rect 559 109 560 111
rect 556 103 560 109
rect 591 128 595 133
rect 600 133 606 142
rect 631 140 633 142
rect 635 140 637 142
rect 631 139 637 140
rect 666 140 668 142
rect 670 140 672 142
rect 600 131 602 133
rect 604 131 606 133
rect 666 135 672 140
rect 688 140 690 142
rect 692 140 694 142
rect 666 133 668 135
rect 670 133 672 135
rect 666 132 672 133
rect 679 134 683 136
rect 679 132 680 134
rect 682 132 683 134
rect 688 135 694 140
rect 688 133 690 135
rect 692 133 694 135
rect 688 132 694 133
rect 720 140 722 142
rect 724 140 726 142
rect 720 135 726 140
rect 742 140 744 142
rect 746 140 748 142
rect 720 133 722 135
rect 724 133 726 135
rect 720 132 726 133
rect 731 134 735 136
rect 731 132 732 134
rect 734 132 735 134
rect 742 135 748 140
rect 777 140 779 142
rect 781 140 783 142
rect 777 139 783 140
rect 818 140 820 142
rect 822 140 824 142
rect 818 139 824 140
rect 742 133 744 135
rect 746 133 748 135
rect 742 132 748 133
rect 799 135 816 136
rect 799 133 801 135
rect 803 133 816 135
rect 799 132 816 133
rect 600 130 606 131
rect 591 126 592 128
rect 594 127 595 128
rect 594 126 608 127
rect 591 123 608 126
rect 542 102 560 103
rect 542 100 544 102
rect 546 100 560 102
rect 542 99 560 100
rect 604 111 608 123
rect 604 109 605 111
rect 607 109 608 111
rect 604 104 608 109
rect 596 100 608 104
rect 596 96 600 100
rect 611 97 612 99
rect 482 93 483 95
rect 485 94 507 95
rect 485 93 503 94
rect 482 92 503 93
rect 505 92 507 94
rect 373 91 398 92
rect 482 91 507 92
rect 512 91 516 93
rect 580 95 600 96
rect 580 93 582 95
rect 584 93 600 95
rect 580 92 600 93
rect 636 128 660 132
rect 679 128 683 132
rect 634 124 640 128
rect 656 127 696 128
rect 656 125 680 127
rect 682 125 696 127
rect 634 114 638 124
rect 644 123 648 125
rect 656 124 696 125
rect 644 121 645 123
rect 647 121 648 123
rect 644 120 648 121
rect 634 112 635 114
rect 637 112 638 114
rect 634 110 638 112
rect 641 116 648 120
rect 641 105 645 116
rect 684 111 688 116
rect 684 109 685 111
rect 687 109 688 111
rect 627 104 645 105
rect 627 102 629 104
rect 631 103 645 104
rect 631 102 656 103
rect 627 101 652 102
rect 641 100 652 101
rect 654 100 656 102
rect 641 99 656 100
rect 661 102 665 104
rect 661 100 662 102
rect 664 100 665 102
rect 661 95 665 100
rect 684 107 688 109
rect 692 113 696 124
rect 692 111 698 113
rect 692 109 695 111
rect 697 109 698 111
rect 692 107 698 109
rect 692 104 696 107
rect 676 100 696 104
rect 676 96 680 100
rect 640 94 662 95
rect 631 91 635 93
rect 640 92 642 94
rect 644 93 662 94
rect 664 93 665 95
rect 644 92 665 93
rect 670 95 680 96
rect 670 93 672 95
rect 674 93 680 95
rect 670 92 680 93
rect 731 128 735 132
rect 754 128 778 132
rect 718 127 758 128
rect 718 125 732 127
rect 734 125 758 127
rect 718 124 758 125
rect 718 113 722 124
rect 766 123 770 125
rect 774 124 780 128
rect 766 121 767 123
rect 769 121 770 123
rect 766 120 770 121
rect 766 116 773 120
rect 716 111 722 113
rect 716 109 717 111
rect 719 109 722 111
rect 716 107 722 109
rect 726 111 730 116
rect 726 109 727 111
rect 729 109 730 111
rect 726 107 730 109
rect 718 104 722 107
rect 718 100 738 104
rect 734 96 738 100
rect 769 105 773 116
rect 776 114 780 124
rect 776 112 777 114
rect 779 112 780 114
rect 776 110 780 112
rect 769 104 787 105
rect 749 102 753 104
rect 769 103 783 104
rect 749 100 750 102
rect 752 100 753 102
rect 734 95 744 96
rect 734 93 740 95
rect 742 93 744 95
rect 734 92 744 93
rect 749 95 753 100
rect 758 102 783 103
rect 785 102 787 104
rect 758 100 760 102
rect 762 101 787 102
rect 762 100 773 101
rect 758 99 773 100
rect 812 128 816 132
rect 812 124 827 128
rect 802 115 808 116
rect 823 111 827 124
rect 830 121 831 132
rect 823 109 824 111
rect 826 109 827 111
rect 823 103 827 109
rect 809 102 827 103
rect 809 100 811 102
rect 813 100 827 102
rect 809 99 827 100
rect 749 93 750 95
rect 752 94 774 95
rect 752 93 770 94
rect 749 92 770 93
rect 772 92 774 94
rect 640 91 665 92
rect 749 91 774 92
rect 779 91 783 93
rect 97 89 98 91
rect 100 89 101 91
rect 245 89 246 91
rect 248 89 249 91
rect 97 86 101 89
rect 153 88 159 89
rect 153 86 155 88
rect 157 86 159 88
rect 187 88 193 89
rect 187 86 189 88
rect 191 86 193 88
rect 245 86 249 89
rect 265 89 271 90
rect 265 87 267 89
rect 269 87 271 89
rect 265 86 271 87
rect 284 89 290 90
rect 284 87 286 89
rect 288 87 290 89
rect 284 86 290 87
rect 364 89 365 91
rect 367 89 368 91
rect 512 89 513 91
rect 515 89 516 91
rect 364 86 368 89
rect 420 88 426 89
rect 420 86 422 88
rect 424 86 426 88
rect 454 88 460 89
rect 454 86 456 88
rect 458 86 460 88
rect 512 86 516 89
rect 532 89 538 90
rect 532 87 534 89
rect 536 87 538 89
rect 532 86 538 87
rect 551 89 557 90
rect 551 87 553 89
rect 555 87 557 89
rect 551 86 557 87
rect 631 89 632 91
rect 634 89 635 91
rect 779 89 780 91
rect 782 89 783 91
rect 631 86 635 89
rect 687 88 693 89
rect 687 86 689 88
rect 691 86 693 88
rect 721 88 727 89
rect 721 86 723 88
rect 725 86 727 88
rect 779 86 783 89
rect 799 89 805 90
rect 799 87 801 89
rect 803 87 805 89
rect 799 86 805 87
rect 818 89 824 90
rect 818 87 820 89
rect 822 87 824 89
rect 818 86 824 87
rect 97 67 101 70
rect 153 68 155 70
rect 157 68 159 70
rect 153 67 159 68
rect 187 68 189 70
rect 191 68 193 70
rect 187 67 193 68
rect 245 67 249 70
rect 97 65 98 67
rect 100 65 101 67
rect 245 65 246 67
rect 248 65 249 67
rect 265 69 271 70
rect 265 67 267 69
rect 269 67 271 69
rect 265 66 271 67
rect 284 69 290 70
rect 284 67 286 69
rect 288 67 290 69
rect 284 66 290 67
rect 364 67 368 70
rect 420 68 422 70
rect 424 68 426 70
rect 420 67 426 68
rect 454 68 456 70
rect 458 68 460 70
rect 454 67 460 68
rect 512 67 516 70
rect 364 65 365 67
rect 367 65 368 67
rect 512 65 513 67
rect 515 65 516 67
rect 532 69 538 70
rect 532 67 534 69
rect 536 67 538 69
rect 532 66 538 67
rect 551 69 557 70
rect 551 67 553 69
rect 555 67 557 69
rect 551 66 557 67
rect 631 67 635 70
rect 687 68 689 70
rect 691 68 693 70
rect 687 67 693 68
rect 721 68 723 70
rect 725 68 727 70
rect 721 67 727 68
rect 779 67 783 70
rect 631 65 632 67
rect 634 65 635 67
rect 779 65 780 67
rect 782 65 783 67
rect 799 69 805 70
rect 799 67 801 69
rect 803 67 805 69
rect 799 66 805 67
rect 818 69 824 70
rect 818 67 820 69
rect 822 67 824 69
rect 818 66 824 67
rect 6 63 26 64
rect 6 61 8 63
rect 10 61 26 63
rect 6 60 26 61
rect 22 56 26 60
rect 46 63 66 64
rect 46 61 48 63
rect 50 61 66 63
rect 46 60 66 61
rect 37 57 38 59
rect 22 52 34 56
rect 30 47 34 52
rect 30 45 31 47
rect 33 45 34 47
rect 30 33 34 45
rect 62 56 66 60
rect 77 57 78 59
rect 62 52 74 56
rect 70 47 74 52
rect 70 45 71 47
rect 73 45 74 47
rect 17 30 34 33
rect 17 28 18 30
rect 20 29 34 30
rect 70 33 74 45
rect 20 28 21 29
rect 6 23 12 24
rect 6 21 8 23
rect 10 21 12 23
rect 6 14 12 21
rect 17 23 21 28
rect 57 30 74 33
rect 57 28 58 30
rect 60 29 74 30
rect 60 28 61 29
rect 17 21 18 23
rect 20 21 21 23
rect 17 19 21 21
rect 26 25 32 26
rect 26 23 28 25
rect 30 23 32 25
rect 26 14 32 23
rect 46 23 52 24
rect 46 21 48 23
rect 50 21 52 23
rect 46 14 52 21
rect 57 23 61 28
rect 97 63 101 65
rect 106 64 131 65
rect 215 64 240 65
rect 106 62 108 64
rect 110 63 131 64
rect 110 62 128 63
rect 106 61 128 62
rect 130 61 131 63
rect 107 56 122 57
rect 107 55 118 56
rect 93 54 118 55
rect 120 54 122 56
rect 93 52 95 54
rect 97 53 122 54
rect 127 56 131 61
rect 136 63 146 64
rect 136 61 138 63
rect 140 61 146 63
rect 136 60 146 61
rect 127 54 128 56
rect 130 54 131 56
rect 97 52 111 53
rect 127 52 131 54
rect 93 51 111 52
rect 100 44 104 46
rect 100 42 101 44
rect 103 42 104 44
rect 100 32 104 42
rect 107 40 111 51
rect 142 56 146 60
rect 142 52 162 56
rect 158 49 162 52
rect 150 47 154 49
rect 150 45 151 47
rect 153 45 154 47
rect 150 40 154 45
rect 158 47 164 49
rect 158 45 161 47
rect 163 45 164 47
rect 158 43 164 45
rect 107 36 114 40
rect 110 35 114 36
rect 110 33 111 35
rect 113 33 114 35
rect 100 28 106 32
rect 110 31 114 33
rect 158 32 162 43
rect 122 31 162 32
rect 122 29 146 31
rect 148 29 162 31
rect 122 28 162 29
rect 57 21 58 23
rect 60 21 61 23
rect 57 19 61 21
rect 66 25 72 26
rect 66 23 68 25
rect 70 23 72 25
rect 102 24 126 28
rect 145 24 149 28
rect 200 63 210 64
rect 200 61 206 63
rect 208 61 210 63
rect 200 60 210 61
rect 215 63 236 64
rect 215 61 216 63
rect 218 62 236 63
rect 238 62 240 64
rect 245 63 249 65
rect 218 61 240 62
rect 200 56 204 60
rect 184 52 204 56
rect 184 49 188 52
rect 182 47 188 49
rect 182 45 183 47
rect 185 45 188 47
rect 182 43 188 45
rect 184 32 188 43
rect 192 47 196 49
rect 215 56 219 61
rect 313 63 333 64
rect 313 61 315 63
rect 317 61 333 63
rect 313 60 333 61
rect 215 54 216 56
rect 218 54 219 56
rect 215 52 219 54
rect 224 56 239 57
rect 224 54 226 56
rect 228 55 239 56
rect 228 54 253 55
rect 224 53 249 54
rect 235 52 249 53
rect 251 52 253 54
rect 235 51 253 52
rect 192 45 193 47
rect 195 45 196 47
rect 192 40 196 45
rect 235 40 239 51
rect 232 36 239 40
rect 242 44 246 46
rect 242 42 243 44
rect 245 42 246 44
rect 232 35 236 36
rect 232 33 233 35
rect 235 33 236 35
rect 184 31 224 32
rect 232 31 236 33
rect 242 32 246 42
rect 275 56 293 57
rect 275 54 277 56
rect 279 54 293 56
rect 275 53 293 54
rect 289 47 293 53
rect 329 56 333 60
rect 344 57 345 59
rect 289 45 290 47
rect 292 45 293 47
rect 268 40 274 41
rect 184 29 198 31
rect 200 29 224 31
rect 184 28 224 29
rect 240 28 246 32
rect 197 24 201 28
rect 220 24 244 28
rect 289 32 293 45
rect 278 28 293 32
rect 278 24 282 28
rect 296 24 297 35
rect 329 52 341 56
rect 337 47 341 52
rect 337 45 338 47
rect 340 45 341 47
rect 337 33 341 45
rect 324 30 341 33
rect 324 28 325 30
rect 327 29 341 30
rect 327 28 328 29
rect 66 14 72 23
rect 132 23 138 24
rect 132 21 134 23
rect 136 21 138 23
rect 97 16 103 17
rect 97 14 99 16
rect 101 14 103 16
rect 132 16 138 21
rect 145 22 146 24
rect 148 22 149 24
rect 145 20 149 22
rect 154 23 160 24
rect 154 21 156 23
rect 158 21 160 23
rect 132 14 134 16
rect 136 14 138 16
rect 154 16 160 21
rect 154 14 156 16
rect 158 14 160 16
rect 186 23 192 24
rect 186 21 188 23
rect 190 21 192 23
rect 186 16 192 21
rect 197 22 198 24
rect 200 22 201 24
rect 197 20 201 22
rect 208 23 214 24
rect 208 21 210 23
rect 212 21 214 23
rect 186 14 188 16
rect 190 14 192 16
rect 208 16 214 21
rect 265 23 282 24
rect 265 21 267 23
rect 269 21 282 23
rect 265 20 282 21
rect 313 23 319 24
rect 313 21 315 23
rect 317 21 319 23
rect 208 14 210 16
rect 212 14 214 16
rect 243 16 249 17
rect 243 14 245 16
rect 247 14 249 16
rect 284 16 290 17
rect 284 14 286 16
rect 288 14 290 16
rect 313 14 319 21
rect 324 23 328 28
rect 364 63 368 65
rect 373 64 398 65
rect 482 64 507 65
rect 373 62 375 64
rect 377 63 398 64
rect 377 62 395 63
rect 373 61 395 62
rect 397 61 398 63
rect 374 56 389 57
rect 374 55 385 56
rect 360 54 385 55
rect 387 54 389 56
rect 360 52 362 54
rect 364 53 389 54
rect 394 56 398 61
rect 403 63 413 64
rect 403 61 405 63
rect 407 61 413 63
rect 403 60 413 61
rect 394 54 395 56
rect 397 54 398 56
rect 364 52 378 53
rect 394 52 398 54
rect 360 51 378 52
rect 367 44 371 46
rect 367 42 368 44
rect 370 42 371 44
rect 367 32 371 42
rect 374 40 378 51
rect 409 56 413 60
rect 409 52 429 56
rect 425 49 429 52
rect 417 47 421 49
rect 417 45 418 47
rect 420 45 421 47
rect 417 40 421 45
rect 425 47 431 49
rect 425 45 428 47
rect 430 45 431 47
rect 425 43 431 45
rect 374 36 381 40
rect 377 35 381 36
rect 377 33 378 35
rect 380 33 381 35
rect 367 28 373 32
rect 377 31 381 33
rect 425 32 429 43
rect 389 31 429 32
rect 389 29 413 31
rect 415 29 429 31
rect 389 28 429 29
rect 324 21 325 23
rect 327 21 328 23
rect 324 19 328 21
rect 333 25 339 26
rect 333 23 335 25
rect 337 23 339 25
rect 369 24 393 28
rect 412 24 416 28
rect 467 63 477 64
rect 467 61 473 63
rect 475 61 477 63
rect 467 60 477 61
rect 482 63 503 64
rect 482 61 483 63
rect 485 62 503 63
rect 505 62 507 64
rect 512 63 516 65
rect 485 61 507 62
rect 467 56 471 60
rect 451 52 471 56
rect 451 49 455 52
rect 449 47 455 49
rect 449 45 450 47
rect 452 45 455 47
rect 449 43 455 45
rect 451 32 455 43
rect 459 47 463 49
rect 482 56 486 61
rect 580 63 600 64
rect 580 61 582 63
rect 584 61 600 63
rect 580 60 600 61
rect 482 54 483 56
rect 485 54 486 56
rect 482 52 486 54
rect 491 56 506 57
rect 491 54 493 56
rect 495 55 506 56
rect 495 54 520 55
rect 491 53 516 54
rect 502 52 516 53
rect 518 52 520 54
rect 502 51 520 52
rect 459 45 460 47
rect 462 45 463 47
rect 459 40 463 45
rect 502 40 506 51
rect 499 36 506 40
rect 509 44 513 46
rect 509 42 510 44
rect 512 42 513 44
rect 499 35 503 36
rect 499 33 500 35
rect 502 33 503 35
rect 451 31 491 32
rect 499 31 503 33
rect 509 32 513 42
rect 542 56 560 57
rect 542 54 544 56
rect 546 54 560 56
rect 542 53 560 54
rect 556 47 560 53
rect 596 56 600 60
rect 611 57 612 59
rect 556 45 557 47
rect 559 45 560 47
rect 535 40 541 41
rect 451 29 465 31
rect 467 29 491 31
rect 451 28 491 29
rect 507 28 513 32
rect 464 24 468 28
rect 487 24 511 28
rect 556 32 560 45
rect 545 28 560 32
rect 545 24 549 28
rect 563 24 564 35
rect 596 52 608 56
rect 604 47 608 52
rect 604 45 605 47
rect 607 45 608 47
rect 604 33 608 45
rect 591 30 608 33
rect 591 28 592 30
rect 594 29 608 30
rect 594 28 595 29
rect 333 14 339 23
rect 399 23 405 24
rect 399 21 401 23
rect 403 21 405 23
rect 364 16 370 17
rect 364 14 366 16
rect 368 14 370 16
rect 399 16 405 21
rect 412 22 413 24
rect 415 22 416 24
rect 412 20 416 22
rect 421 23 427 24
rect 421 21 423 23
rect 425 21 427 23
rect 399 14 401 16
rect 403 14 405 16
rect 421 16 427 21
rect 421 14 423 16
rect 425 14 427 16
rect 453 23 459 24
rect 453 21 455 23
rect 457 21 459 23
rect 453 16 459 21
rect 464 22 465 24
rect 467 22 468 24
rect 464 20 468 22
rect 475 23 481 24
rect 475 21 477 23
rect 479 21 481 23
rect 453 14 455 16
rect 457 14 459 16
rect 475 16 481 21
rect 532 23 549 24
rect 532 21 534 23
rect 536 21 549 23
rect 532 20 549 21
rect 580 23 586 24
rect 580 21 582 23
rect 584 21 586 23
rect 475 14 477 16
rect 479 14 481 16
rect 510 16 516 17
rect 510 14 512 16
rect 514 14 516 16
rect 551 16 557 17
rect 551 14 553 16
rect 555 14 557 16
rect 580 14 586 21
rect 591 23 595 28
rect 631 63 635 65
rect 640 64 665 65
rect 749 64 774 65
rect 640 62 642 64
rect 644 63 665 64
rect 644 62 662 63
rect 640 61 662 62
rect 664 61 665 63
rect 641 56 656 57
rect 641 55 652 56
rect 627 54 652 55
rect 654 54 656 56
rect 627 52 629 54
rect 631 53 656 54
rect 661 56 665 61
rect 670 63 680 64
rect 670 61 672 63
rect 674 61 680 63
rect 670 60 680 61
rect 661 54 662 56
rect 664 54 665 56
rect 631 52 645 53
rect 661 52 665 54
rect 627 51 645 52
rect 634 44 638 46
rect 634 42 635 44
rect 637 42 638 44
rect 634 32 638 42
rect 641 40 645 51
rect 676 56 680 60
rect 676 52 696 56
rect 692 49 696 52
rect 684 47 688 49
rect 684 45 685 47
rect 687 45 688 47
rect 684 40 688 45
rect 692 47 698 49
rect 692 45 695 47
rect 697 45 698 47
rect 692 43 698 45
rect 641 36 648 40
rect 644 35 648 36
rect 644 33 645 35
rect 647 33 648 35
rect 634 28 640 32
rect 644 31 648 33
rect 692 32 696 43
rect 656 31 696 32
rect 656 29 680 31
rect 682 29 696 31
rect 656 28 696 29
rect 591 21 592 23
rect 594 21 595 23
rect 591 19 595 21
rect 600 25 606 26
rect 600 23 602 25
rect 604 23 606 25
rect 636 24 660 28
rect 679 24 683 28
rect 734 63 744 64
rect 734 61 740 63
rect 742 61 744 63
rect 734 60 744 61
rect 749 63 770 64
rect 749 61 750 63
rect 752 62 770 63
rect 772 62 774 64
rect 779 63 783 65
rect 752 61 774 62
rect 734 56 738 60
rect 718 52 738 56
rect 718 49 722 52
rect 716 47 722 49
rect 716 45 717 47
rect 719 45 722 47
rect 716 43 722 45
rect 718 32 722 43
rect 726 47 730 49
rect 749 56 753 61
rect 749 54 750 56
rect 752 54 753 56
rect 749 52 753 54
rect 758 56 773 57
rect 758 54 760 56
rect 762 55 773 56
rect 762 54 787 55
rect 758 53 783 54
rect 769 52 783 53
rect 785 52 787 54
rect 769 51 787 52
rect 726 45 727 47
rect 729 45 730 47
rect 726 40 730 45
rect 769 40 773 51
rect 766 36 773 40
rect 776 44 780 46
rect 776 42 777 44
rect 779 42 780 44
rect 766 35 770 36
rect 766 33 767 35
rect 769 33 770 35
rect 718 31 758 32
rect 766 31 770 33
rect 776 32 780 42
rect 809 56 827 57
rect 809 54 811 56
rect 813 54 827 56
rect 809 53 827 54
rect 823 47 827 53
rect 823 45 824 47
rect 826 45 827 47
rect 802 40 808 41
rect 718 29 732 31
rect 734 29 758 31
rect 718 28 758 29
rect 774 28 780 32
rect 731 24 735 28
rect 754 24 778 28
rect 823 32 827 45
rect 812 28 827 32
rect 812 24 816 28
rect 830 24 831 35
rect 600 14 606 23
rect 666 23 672 24
rect 666 21 668 23
rect 670 21 672 23
rect 631 16 637 17
rect 631 14 633 16
rect 635 14 637 16
rect 666 16 672 21
rect 679 22 680 24
rect 682 22 683 24
rect 679 20 683 22
rect 688 23 694 24
rect 688 21 690 23
rect 692 21 694 23
rect 666 14 668 16
rect 670 14 672 16
rect 688 16 694 21
rect 688 14 690 16
rect 692 14 694 16
rect 720 23 726 24
rect 720 21 722 23
rect 724 21 726 23
rect 720 16 726 21
rect 731 22 732 24
rect 734 22 735 24
rect 731 20 735 22
rect 742 23 748 24
rect 742 21 744 23
rect 746 21 748 23
rect 720 14 722 16
rect 724 14 726 16
rect 742 16 748 21
rect 799 23 816 24
rect 799 21 801 23
rect 803 21 816 23
rect 799 20 816 21
rect 742 14 744 16
rect 746 14 748 16
rect 777 16 783 17
rect 777 14 779 16
rect 781 14 783 16
rect 818 16 824 17
rect 818 14 820 16
rect 822 14 824 16
rect 443 -4 444 -2
rect 446 -4 447 -2
rect 443 -9 447 -4
rect 499 -4 501 -2
rect 503 -4 505 -2
rect 499 -5 505 -4
rect 534 -4 536 -2
rect 538 -4 540 -2
rect 443 -11 444 -9
rect 446 -11 447 -9
rect 443 -13 447 -11
rect 451 -8 484 -7
rect 451 -10 480 -8
rect 482 -10 484 -8
rect 451 -11 484 -10
rect 534 -9 540 -4
rect 556 -4 558 -2
rect 560 -4 562 -2
rect 534 -11 536 -9
rect 538 -11 540 -9
rect 451 -22 455 -11
rect 534 -12 540 -11
rect 547 -10 551 -8
rect 547 -12 548 -10
rect 550 -12 551 -10
rect 556 -9 562 -4
rect 556 -11 558 -9
rect 560 -11 562 -9
rect 556 -12 562 -11
rect 588 -4 590 -2
rect 592 -4 594 -2
rect 588 -9 594 -4
rect 610 -4 612 -2
rect 614 -4 616 -2
rect 588 -11 590 -9
rect 592 -11 594 -9
rect 588 -12 594 -11
rect 599 -10 603 -8
rect 599 -12 600 -10
rect 602 -12 603 -10
rect 610 -9 616 -4
rect 645 -4 647 -2
rect 649 -4 651 -2
rect 645 -5 651 -4
rect 686 -4 688 -2
rect 690 -4 692 -2
rect 686 -5 692 -4
rect 721 -4 722 -2
rect 724 -4 725 -2
rect 721 -6 725 -4
rect 754 -4 756 -2
rect 758 -4 760 -2
rect 754 -5 760 -4
rect 785 -4 786 -2
rect 788 -4 789 -2
rect 785 -6 789 -4
rect 818 -4 820 -2
rect 822 -4 824 -2
rect 818 -5 824 -4
rect 610 -11 612 -9
rect 614 -11 616 -9
rect 610 -12 616 -11
rect 667 -9 684 -8
rect 667 -11 669 -9
rect 671 -11 684 -9
rect 667 -12 684 -11
rect 432 -23 455 -22
rect 432 -25 434 -23
rect 436 -25 455 -23
rect 432 -26 455 -25
rect 432 -32 436 -26
rect 425 -36 436 -32
rect 425 -42 429 -36
rect 451 -32 455 -26
rect 459 -16 463 -14
rect 459 -18 460 -16
rect 462 -18 463 -16
rect 459 -23 463 -18
rect 459 -25 460 -23
rect 462 -24 463 -23
rect 462 -25 475 -24
rect 459 -28 475 -25
rect 471 -30 475 -28
rect 471 -32 476 -30
rect 451 -33 467 -32
rect 451 -35 463 -33
rect 465 -35 467 -33
rect 451 -36 467 -35
rect 471 -34 473 -32
rect 475 -34 476 -32
rect 471 -36 476 -34
rect 425 -44 426 -42
rect 428 -44 429 -42
rect 425 -46 429 -44
rect 471 -40 475 -36
rect 451 -44 475 -40
rect 451 -47 455 -44
rect 451 -49 452 -47
rect 454 -49 455 -47
rect 438 -50 444 -49
rect 438 -52 440 -50
rect 442 -52 444 -50
rect 451 -51 455 -49
rect 504 -16 528 -12
rect 547 -16 551 -12
rect 502 -20 508 -16
rect 524 -17 564 -16
rect 524 -19 548 -17
rect 550 -19 564 -17
rect 502 -30 506 -20
rect 512 -21 516 -19
rect 524 -20 564 -19
rect 512 -23 513 -21
rect 515 -23 516 -21
rect 512 -24 516 -23
rect 502 -32 503 -30
rect 505 -32 506 -30
rect 502 -34 506 -32
rect 509 -28 516 -24
rect 509 -39 513 -28
rect 552 -33 556 -28
rect 552 -35 553 -33
rect 555 -35 556 -33
rect 495 -40 513 -39
rect 495 -42 497 -40
rect 499 -41 513 -40
rect 499 -42 524 -41
rect 495 -43 520 -42
rect 509 -44 520 -43
rect 522 -44 524 -42
rect 509 -45 524 -44
rect 529 -42 533 -40
rect 529 -44 530 -42
rect 532 -44 533 -42
rect 529 -49 533 -44
rect 552 -37 556 -35
rect 560 -31 564 -20
rect 560 -33 566 -31
rect 560 -35 563 -33
rect 565 -35 566 -33
rect 560 -37 566 -35
rect 560 -40 564 -37
rect 544 -44 564 -40
rect 544 -48 548 -44
rect 508 -50 530 -49
rect 438 -58 444 -52
rect 499 -53 503 -51
rect 508 -52 510 -50
rect 512 -51 530 -50
rect 532 -51 533 -49
rect 512 -52 533 -51
rect 538 -49 548 -48
rect 538 -51 540 -49
rect 542 -51 548 -49
rect 538 -52 548 -51
rect 599 -16 603 -12
rect 622 -16 646 -12
rect 586 -17 626 -16
rect 586 -19 600 -17
rect 602 -19 626 -17
rect 586 -20 626 -19
rect 586 -31 590 -20
rect 634 -21 638 -19
rect 642 -20 648 -16
rect 634 -23 635 -21
rect 637 -23 638 -21
rect 634 -24 638 -23
rect 634 -28 641 -24
rect 584 -33 590 -31
rect 584 -35 585 -33
rect 587 -35 590 -33
rect 584 -37 590 -35
rect 594 -33 598 -28
rect 594 -35 595 -33
rect 597 -35 598 -33
rect 594 -37 598 -35
rect 586 -40 590 -37
rect 586 -44 606 -40
rect 602 -48 606 -44
rect 637 -39 641 -28
rect 644 -30 648 -20
rect 644 -32 645 -30
rect 647 -32 648 -30
rect 644 -34 648 -32
rect 637 -40 655 -39
rect 617 -42 621 -40
rect 637 -41 651 -40
rect 617 -44 618 -42
rect 620 -44 621 -42
rect 602 -49 612 -48
rect 602 -51 608 -49
rect 610 -51 612 -49
rect 602 -52 612 -51
rect 617 -49 621 -44
rect 626 -42 651 -41
rect 653 -42 655 -40
rect 626 -44 628 -42
rect 630 -43 655 -42
rect 630 -44 641 -43
rect 626 -45 641 -44
rect 680 -16 684 -12
rect 680 -20 695 -16
rect 670 -29 676 -28
rect 691 -33 695 -20
rect 698 -23 699 -12
rect 737 -12 750 -11
rect 737 -14 739 -12
rect 741 -14 750 -12
rect 737 -15 750 -14
rect 746 -19 762 -15
rect 691 -35 692 -33
rect 694 -35 695 -33
rect 691 -41 695 -35
rect 734 -23 738 -21
rect 677 -42 695 -41
rect 677 -44 679 -42
rect 681 -44 695 -42
rect 677 -45 695 -44
rect 710 -24 735 -23
rect 710 -26 712 -24
rect 714 -25 735 -24
rect 737 -25 738 -23
rect 714 -26 738 -25
rect 710 -27 738 -26
rect 710 -47 714 -27
rect 734 -37 738 -27
rect 754 -32 755 -26
rect 758 -36 762 -19
rect 734 -39 745 -37
rect 734 -41 742 -39
rect 744 -41 745 -39
rect 758 -38 763 -36
rect 758 -40 760 -38
rect 762 -40 763 -38
rect 734 -43 745 -41
rect 748 -42 763 -40
rect 748 -44 762 -42
rect 710 -48 716 -47
rect 617 -51 618 -49
rect 620 -50 642 -49
rect 620 -51 638 -50
rect 617 -52 638 -51
rect 640 -52 642 -50
rect 710 -50 712 -48
rect 714 -50 716 -48
rect 710 -51 716 -50
rect 720 -48 726 -47
rect 720 -50 722 -48
rect 724 -50 726 -48
rect 748 -49 752 -44
rect 801 -12 814 -11
rect 801 -14 803 -12
rect 805 -14 814 -12
rect 801 -15 814 -14
rect 810 -19 826 -15
rect 798 -23 802 -21
rect 508 -53 533 -52
rect 617 -53 642 -52
rect 647 -53 651 -51
rect 499 -55 500 -53
rect 502 -55 503 -53
rect 647 -55 648 -53
rect 650 -55 651 -53
rect 499 -58 503 -55
rect 555 -56 561 -55
rect 555 -58 557 -56
rect 559 -58 561 -56
rect 589 -56 595 -55
rect 589 -58 591 -56
rect 593 -58 595 -56
rect 647 -58 651 -55
rect 667 -55 673 -54
rect 667 -57 669 -55
rect 671 -57 673 -55
rect 667 -58 673 -57
rect 686 -55 692 -54
rect 686 -57 688 -55
rect 690 -57 692 -55
rect 686 -58 692 -57
rect 720 -58 726 -50
rect 737 -50 752 -49
rect 737 -52 739 -50
rect 741 -52 752 -50
rect 737 -53 752 -52
rect 755 -50 759 -48
rect 755 -52 756 -50
rect 758 -52 759 -50
rect 755 -58 759 -52
rect 774 -24 799 -23
rect 774 -26 776 -24
rect 778 -25 799 -24
rect 801 -25 802 -23
rect 778 -26 802 -25
rect 774 -27 802 -26
rect 774 -47 778 -27
rect 798 -37 802 -27
rect 818 -32 819 -26
rect 822 -36 826 -19
rect 798 -39 809 -37
rect 798 -41 806 -39
rect 808 -41 809 -39
rect 822 -38 827 -36
rect 822 -40 824 -38
rect 826 -40 827 -38
rect 798 -43 809 -41
rect 812 -42 827 -40
rect 812 -44 826 -42
rect 774 -48 780 -47
rect 774 -50 776 -48
rect 778 -50 780 -48
rect 774 -51 780 -50
rect 784 -48 790 -47
rect 784 -50 786 -48
rect 788 -50 790 -48
rect 812 -49 816 -44
rect 784 -58 790 -50
rect 801 -50 816 -49
rect 801 -52 803 -50
rect 805 -52 816 -50
rect 801 -53 816 -52
rect 819 -50 823 -48
rect 819 -52 820 -50
rect 822 -52 823 -50
rect 819 -58 823 -52
rect 438 -80 444 -74
rect 499 -77 503 -74
rect 555 -76 557 -74
rect 559 -76 561 -74
rect 555 -77 561 -76
rect 589 -76 591 -74
rect 593 -76 595 -74
rect 589 -77 595 -76
rect 647 -77 651 -74
rect 499 -79 500 -77
rect 502 -79 503 -77
rect 647 -79 648 -77
rect 650 -79 651 -77
rect 667 -75 673 -74
rect 667 -77 669 -75
rect 671 -77 673 -75
rect 667 -78 673 -77
rect 686 -75 692 -74
rect 686 -77 688 -75
rect 690 -77 692 -75
rect 686 -78 692 -77
rect 438 -82 440 -80
rect 442 -82 444 -80
rect 438 -83 444 -82
rect 451 -83 455 -81
rect 451 -85 452 -83
rect 454 -85 455 -83
rect 425 -88 429 -86
rect 425 -90 426 -88
rect 428 -90 429 -88
rect 425 -96 429 -90
rect 451 -88 455 -85
rect 451 -92 475 -88
rect 425 -100 436 -96
rect 432 -106 436 -100
rect 471 -96 475 -92
rect 451 -97 467 -96
rect 451 -99 463 -97
rect 465 -99 467 -97
rect 451 -100 467 -99
rect 471 -98 476 -96
rect 471 -100 473 -98
rect 475 -100 476 -98
rect 451 -106 455 -100
rect 471 -102 476 -100
rect 471 -104 475 -102
rect 432 -107 455 -106
rect 432 -109 434 -107
rect 436 -109 455 -107
rect 432 -110 455 -109
rect 443 -121 447 -119
rect 443 -123 444 -121
rect 446 -123 447 -121
rect 443 -128 447 -123
rect 451 -121 455 -110
rect 459 -107 475 -104
rect 459 -109 460 -107
rect 462 -108 475 -107
rect 462 -109 463 -108
rect 459 -114 463 -109
rect 459 -116 460 -114
rect 462 -116 463 -114
rect 459 -118 463 -116
rect 499 -81 503 -79
rect 508 -80 533 -79
rect 617 -80 642 -79
rect 508 -82 510 -80
rect 512 -81 533 -80
rect 512 -82 530 -81
rect 508 -83 530 -82
rect 532 -83 533 -81
rect 509 -88 524 -87
rect 509 -89 520 -88
rect 495 -90 520 -89
rect 522 -90 524 -88
rect 495 -92 497 -90
rect 499 -91 524 -90
rect 529 -88 533 -83
rect 538 -81 548 -80
rect 538 -83 540 -81
rect 542 -83 548 -81
rect 538 -84 548 -83
rect 529 -90 530 -88
rect 532 -90 533 -88
rect 499 -92 513 -91
rect 529 -92 533 -90
rect 495 -93 513 -92
rect 502 -100 506 -98
rect 502 -102 503 -100
rect 505 -102 506 -100
rect 502 -112 506 -102
rect 509 -104 513 -93
rect 544 -88 548 -84
rect 544 -92 564 -88
rect 560 -95 564 -92
rect 552 -97 556 -95
rect 552 -99 553 -97
rect 555 -99 556 -97
rect 552 -104 556 -99
rect 560 -97 566 -95
rect 560 -99 563 -97
rect 565 -99 566 -97
rect 560 -101 566 -99
rect 509 -108 516 -104
rect 512 -109 516 -108
rect 512 -111 513 -109
rect 515 -111 516 -109
rect 502 -116 508 -112
rect 512 -113 516 -111
rect 560 -112 564 -101
rect 524 -113 564 -112
rect 524 -115 548 -113
rect 550 -115 564 -113
rect 524 -116 564 -115
rect 504 -120 528 -116
rect 547 -120 551 -116
rect 602 -81 612 -80
rect 602 -83 608 -81
rect 610 -83 612 -81
rect 602 -84 612 -83
rect 617 -81 638 -80
rect 617 -83 618 -81
rect 620 -82 638 -81
rect 640 -82 642 -80
rect 647 -81 651 -79
rect 620 -83 642 -82
rect 602 -88 606 -84
rect 586 -92 606 -88
rect 586 -95 590 -92
rect 584 -97 590 -95
rect 584 -99 585 -97
rect 587 -99 590 -97
rect 584 -101 590 -99
rect 586 -112 590 -101
rect 594 -97 598 -95
rect 617 -88 621 -83
rect 710 -82 716 -81
rect 710 -84 712 -82
rect 714 -84 716 -82
rect 617 -90 618 -88
rect 620 -90 621 -88
rect 617 -92 621 -90
rect 626 -88 641 -87
rect 626 -90 628 -88
rect 630 -89 641 -88
rect 630 -90 655 -89
rect 626 -91 651 -90
rect 637 -92 651 -91
rect 653 -92 655 -90
rect 637 -93 655 -92
rect 594 -99 595 -97
rect 597 -99 598 -97
rect 594 -104 598 -99
rect 637 -104 641 -93
rect 634 -108 641 -104
rect 644 -100 648 -98
rect 644 -102 645 -100
rect 647 -102 648 -100
rect 634 -109 638 -108
rect 634 -111 635 -109
rect 637 -111 638 -109
rect 586 -113 626 -112
rect 634 -113 638 -111
rect 644 -112 648 -102
rect 710 -85 716 -84
rect 720 -82 726 -74
rect 720 -84 722 -82
rect 724 -84 726 -82
rect 737 -80 752 -79
rect 737 -82 739 -80
rect 741 -82 752 -80
rect 737 -83 752 -82
rect 720 -85 726 -84
rect 677 -88 695 -87
rect 677 -90 679 -88
rect 681 -90 695 -88
rect 677 -91 695 -90
rect 691 -97 695 -91
rect 691 -99 692 -97
rect 694 -99 695 -97
rect 670 -104 676 -103
rect 586 -115 600 -113
rect 602 -115 626 -113
rect 586 -116 626 -115
rect 642 -116 648 -112
rect 599 -120 603 -116
rect 622 -120 646 -116
rect 691 -112 695 -99
rect 680 -116 695 -112
rect 680 -120 684 -116
rect 698 -120 699 -109
rect 710 -105 714 -85
rect 748 -88 752 -83
rect 755 -80 759 -74
rect 755 -82 756 -80
rect 758 -82 759 -80
rect 755 -84 759 -82
rect 734 -91 745 -89
rect 734 -93 742 -91
rect 744 -93 745 -91
rect 748 -90 762 -88
rect 748 -92 763 -90
rect 734 -95 745 -93
rect 758 -94 760 -92
rect 762 -94 763 -92
rect 734 -105 738 -95
rect 758 -96 763 -94
rect 710 -106 738 -105
rect 710 -108 712 -106
rect 714 -107 738 -106
rect 714 -108 735 -107
rect 710 -109 735 -108
rect 737 -109 738 -107
rect 754 -106 755 -100
rect 734 -111 738 -109
rect 534 -121 540 -120
rect 451 -122 484 -121
rect 451 -124 480 -122
rect 482 -124 484 -122
rect 451 -125 484 -124
rect 534 -123 536 -121
rect 538 -123 540 -121
rect 443 -130 444 -128
rect 446 -130 447 -128
rect 499 -128 505 -127
rect 499 -130 501 -128
rect 503 -130 505 -128
rect 534 -128 540 -123
rect 547 -122 548 -120
rect 550 -122 551 -120
rect 547 -124 551 -122
rect 556 -121 562 -120
rect 556 -123 558 -121
rect 560 -123 562 -121
rect 534 -130 536 -128
rect 538 -130 540 -128
rect 556 -128 562 -123
rect 556 -130 558 -128
rect 560 -130 562 -128
rect 588 -121 594 -120
rect 588 -123 590 -121
rect 592 -123 594 -121
rect 588 -128 594 -123
rect 599 -122 600 -120
rect 602 -122 603 -120
rect 599 -124 603 -122
rect 610 -121 616 -120
rect 610 -123 612 -121
rect 614 -123 616 -121
rect 588 -130 590 -128
rect 592 -130 594 -128
rect 610 -128 616 -123
rect 667 -121 684 -120
rect 667 -123 669 -121
rect 671 -123 684 -121
rect 667 -124 684 -123
rect 758 -113 762 -96
rect 746 -117 762 -113
rect 737 -118 750 -117
rect 737 -120 739 -118
rect 741 -120 750 -118
rect 774 -82 780 -81
rect 774 -84 776 -82
rect 778 -84 780 -82
rect 774 -85 780 -84
rect 784 -82 790 -74
rect 784 -84 786 -82
rect 788 -84 790 -82
rect 801 -80 816 -79
rect 801 -82 803 -80
rect 805 -82 816 -80
rect 801 -83 816 -82
rect 784 -85 790 -84
rect 774 -105 778 -85
rect 812 -88 816 -83
rect 819 -80 823 -74
rect 819 -82 820 -80
rect 822 -82 823 -80
rect 819 -84 823 -82
rect 798 -91 809 -89
rect 798 -93 806 -91
rect 808 -93 809 -91
rect 812 -90 826 -88
rect 812 -92 827 -90
rect 798 -95 809 -93
rect 822 -94 824 -92
rect 826 -94 827 -92
rect 798 -105 802 -95
rect 822 -96 827 -94
rect 774 -106 802 -105
rect 774 -108 776 -106
rect 778 -107 802 -106
rect 778 -108 799 -107
rect 774 -109 799 -108
rect 801 -109 802 -107
rect 818 -106 819 -100
rect 798 -111 802 -109
rect 737 -121 750 -120
rect 822 -113 826 -96
rect 810 -117 826 -113
rect 801 -118 814 -117
rect 801 -120 803 -118
rect 805 -120 814 -118
rect 801 -121 814 -120
rect 610 -130 612 -128
rect 614 -130 616 -128
rect 645 -128 651 -127
rect 645 -130 647 -128
rect 649 -130 651 -128
rect 686 -128 692 -127
rect 686 -130 688 -128
rect 690 -130 692 -128
rect 721 -128 725 -126
rect 721 -130 722 -128
rect 724 -130 725 -128
rect 754 -128 760 -127
rect 754 -130 756 -128
rect 758 -130 760 -128
rect 785 -128 789 -126
rect 785 -130 786 -128
rect 788 -130 789 -128
rect 818 -128 824 -127
rect 818 -130 820 -128
rect 822 -130 824 -128
rect 443 -148 444 -146
rect 446 -148 447 -146
rect 443 -153 447 -148
rect 499 -148 501 -146
rect 503 -148 505 -146
rect 499 -149 505 -148
rect 534 -148 536 -146
rect 538 -148 540 -146
rect 443 -155 444 -153
rect 446 -155 447 -153
rect 443 -157 447 -155
rect 451 -152 484 -151
rect 451 -154 480 -152
rect 482 -154 484 -152
rect 451 -155 484 -154
rect 534 -153 540 -148
rect 556 -148 558 -146
rect 560 -148 562 -146
rect 534 -155 536 -153
rect 538 -155 540 -153
rect 451 -166 455 -155
rect 534 -156 540 -155
rect 547 -154 551 -152
rect 547 -156 548 -154
rect 550 -156 551 -154
rect 556 -153 562 -148
rect 556 -155 558 -153
rect 560 -155 562 -153
rect 556 -156 562 -155
rect 588 -148 590 -146
rect 592 -148 594 -146
rect 588 -153 594 -148
rect 610 -148 612 -146
rect 614 -148 616 -146
rect 588 -155 590 -153
rect 592 -155 594 -153
rect 588 -156 594 -155
rect 599 -154 603 -152
rect 599 -156 600 -154
rect 602 -156 603 -154
rect 610 -153 616 -148
rect 645 -148 647 -146
rect 649 -148 651 -146
rect 645 -149 651 -148
rect 686 -148 688 -146
rect 690 -148 692 -146
rect 686 -149 692 -148
rect 721 -148 722 -146
rect 724 -148 725 -146
rect 721 -150 725 -148
rect 754 -148 756 -146
rect 758 -148 760 -146
rect 754 -149 760 -148
rect 785 -148 786 -146
rect 788 -148 789 -146
rect 785 -150 789 -148
rect 818 -148 820 -146
rect 822 -148 824 -146
rect 818 -149 824 -148
rect 610 -155 612 -153
rect 614 -155 616 -153
rect 610 -156 616 -155
rect 667 -153 684 -152
rect 667 -155 669 -153
rect 671 -155 684 -153
rect 667 -156 684 -155
rect 432 -167 455 -166
rect 432 -169 434 -167
rect 436 -169 455 -167
rect 432 -170 455 -169
rect 432 -176 436 -170
rect 425 -180 436 -176
rect 425 -186 429 -180
rect 451 -176 455 -170
rect 459 -160 463 -158
rect 459 -162 460 -160
rect 462 -162 463 -160
rect 459 -167 463 -162
rect 459 -169 460 -167
rect 462 -168 463 -167
rect 462 -169 475 -168
rect 459 -172 475 -169
rect 471 -174 475 -172
rect 471 -176 476 -174
rect 451 -177 467 -176
rect 451 -179 463 -177
rect 465 -179 467 -177
rect 451 -180 467 -179
rect 471 -178 473 -176
rect 475 -178 476 -176
rect 471 -180 476 -178
rect 425 -188 426 -186
rect 428 -188 429 -186
rect 425 -190 429 -188
rect 471 -184 475 -180
rect 451 -188 475 -184
rect 451 -191 455 -188
rect 451 -193 452 -191
rect 454 -193 455 -191
rect 438 -194 444 -193
rect 438 -196 440 -194
rect 442 -196 444 -194
rect 451 -195 455 -193
rect 504 -160 528 -156
rect 547 -160 551 -156
rect 502 -164 508 -160
rect 524 -161 564 -160
rect 524 -163 548 -161
rect 550 -163 564 -161
rect 502 -174 506 -164
rect 512 -165 516 -163
rect 524 -164 564 -163
rect 512 -167 513 -165
rect 515 -167 516 -165
rect 512 -168 516 -167
rect 502 -176 503 -174
rect 505 -176 506 -174
rect 502 -178 506 -176
rect 509 -172 516 -168
rect 509 -183 513 -172
rect 552 -177 556 -172
rect 552 -179 553 -177
rect 555 -179 556 -177
rect 495 -184 513 -183
rect 495 -186 497 -184
rect 499 -185 513 -184
rect 499 -186 524 -185
rect 495 -187 520 -186
rect 509 -188 520 -187
rect 522 -188 524 -186
rect 509 -189 524 -188
rect 529 -186 533 -184
rect 529 -188 530 -186
rect 532 -188 533 -186
rect 529 -193 533 -188
rect 552 -181 556 -179
rect 560 -175 564 -164
rect 560 -177 566 -175
rect 560 -179 563 -177
rect 565 -179 566 -177
rect 560 -181 566 -179
rect 560 -184 564 -181
rect 544 -188 564 -184
rect 544 -192 548 -188
rect 508 -194 530 -193
rect 438 -202 444 -196
rect 499 -197 503 -195
rect 508 -196 510 -194
rect 512 -195 530 -194
rect 532 -195 533 -193
rect 512 -196 533 -195
rect 538 -193 548 -192
rect 538 -195 540 -193
rect 542 -195 548 -193
rect 538 -196 548 -195
rect 599 -160 603 -156
rect 622 -160 646 -156
rect 586 -161 626 -160
rect 586 -163 600 -161
rect 602 -163 626 -161
rect 586 -164 626 -163
rect 586 -175 590 -164
rect 634 -165 638 -163
rect 642 -164 648 -160
rect 634 -167 635 -165
rect 637 -167 638 -165
rect 634 -168 638 -167
rect 634 -172 641 -168
rect 584 -177 590 -175
rect 584 -179 585 -177
rect 587 -179 590 -177
rect 584 -181 590 -179
rect 594 -177 598 -172
rect 594 -179 595 -177
rect 597 -179 598 -177
rect 594 -181 598 -179
rect 586 -184 590 -181
rect 586 -188 606 -184
rect 602 -192 606 -188
rect 637 -183 641 -172
rect 644 -174 648 -164
rect 644 -176 645 -174
rect 647 -176 648 -174
rect 644 -178 648 -176
rect 637 -184 655 -183
rect 617 -186 621 -184
rect 637 -185 651 -184
rect 617 -188 618 -186
rect 620 -188 621 -186
rect 602 -193 612 -192
rect 602 -195 608 -193
rect 610 -195 612 -193
rect 602 -196 612 -195
rect 617 -193 621 -188
rect 626 -186 651 -185
rect 653 -186 655 -184
rect 626 -188 628 -186
rect 630 -187 655 -186
rect 630 -188 641 -187
rect 626 -189 641 -188
rect 680 -160 684 -156
rect 680 -164 695 -160
rect 670 -173 676 -172
rect 691 -177 695 -164
rect 698 -167 699 -156
rect 737 -156 750 -155
rect 737 -158 739 -156
rect 741 -158 750 -156
rect 737 -159 750 -158
rect 746 -163 762 -159
rect 691 -179 692 -177
rect 694 -179 695 -177
rect 691 -185 695 -179
rect 734 -167 738 -165
rect 677 -186 695 -185
rect 677 -188 679 -186
rect 681 -188 695 -186
rect 677 -189 695 -188
rect 710 -168 735 -167
rect 710 -170 712 -168
rect 714 -169 735 -168
rect 737 -169 738 -167
rect 714 -170 738 -169
rect 710 -171 738 -170
rect 710 -191 714 -171
rect 734 -181 738 -171
rect 754 -176 755 -170
rect 758 -180 762 -163
rect 801 -156 814 -155
rect 801 -158 803 -156
rect 805 -158 814 -156
rect 801 -159 814 -158
rect 810 -163 826 -159
rect 798 -167 802 -165
rect 734 -183 745 -181
rect 734 -185 742 -183
rect 744 -185 745 -183
rect 758 -182 763 -180
rect 758 -184 760 -182
rect 762 -184 763 -182
rect 734 -187 745 -185
rect 748 -186 763 -184
rect 748 -188 762 -186
rect 617 -195 618 -193
rect 620 -194 642 -193
rect 620 -195 638 -194
rect 617 -196 638 -195
rect 640 -196 642 -194
rect 710 -192 716 -191
rect 710 -194 712 -192
rect 714 -194 716 -192
rect 710 -195 716 -194
rect 720 -192 726 -191
rect 720 -194 722 -192
rect 724 -194 726 -192
rect 748 -193 752 -188
rect 508 -197 533 -196
rect 617 -197 642 -196
rect 647 -197 651 -195
rect 499 -199 500 -197
rect 502 -199 503 -197
rect 647 -199 648 -197
rect 650 -199 651 -197
rect 499 -202 503 -199
rect 555 -200 561 -199
rect 555 -202 557 -200
rect 559 -202 561 -200
rect 589 -200 595 -199
rect 589 -202 591 -200
rect 593 -202 595 -200
rect 647 -202 651 -199
rect 667 -199 673 -198
rect 667 -201 669 -199
rect 671 -201 673 -199
rect 667 -202 673 -201
rect 686 -199 692 -198
rect 686 -201 688 -199
rect 690 -201 692 -199
rect 686 -202 692 -201
rect 720 -202 726 -194
rect 737 -194 752 -193
rect 737 -196 739 -194
rect 741 -196 752 -194
rect 737 -197 752 -196
rect 755 -194 759 -192
rect 755 -196 756 -194
rect 758 -196 759 -194
rect 774 -168 799 -167
rect 774 -170 776 -168
rect 778 -169 799 -168
rect 801 -169 802 -167
rect 778 -170 802 -169
rect 774 -171 802 -170
rect 774 -191 778 -171
rect 798 -181 802 -171
rect 818 -176 819 -170
rect 822 -180 826 -163
rect 798 -183 809 -181
rect 798 -185 806 -183
rect 808 -185 809 -183
rect 822 -182 827 -180
rect 822 -184 824 -182
rect 826 -184 827 -182
rect 798 -187 809 -185
rect 812 -186 827 -184
rect 812 -188 826 -186
rect 774 -192 780 -191
rect 774 -194 776 -192
rect 778 -194 780 -192
rect 774 -195 780 -194
rect 784 -192 790 -191
rect 784 -194 786 -192
rect 788 -194 790 -192
rect 812 -193 816 -188
rect 755 -202 759 -196
rect 784 -202 790 -194
rect 801 -194 816 -193
rect 801 -196 803 -194
rect 805 -196 816 -194
rect 801 -197 816 -196
rect 819 -194 823 -192
rect 819 -196 820 -194
rect 822 -196 823 -194
rect 819 -202 823 -196
rect 438 -224 444 -218
rect 499 -221 503 -218
rect 555 -220 557 -218
rect 559 -220 561 -218
rect 555 -221 561 -220
rect 589 -220 591 -218
rect 593 -220 595 -218
rect 589 -221 595 -220
rect 647 -221 651 -218
rect 499 -223 500 -221
rect 502 -223 503 -221
rect 647 -223 648 -221
rect 650 -223 651 -221
rect 667 -219 673 -218
rect 667 -221 669 -219
rect 671 -221 673 -219
rect 667 -222 673 -221
rect 686 -219 692 -218
rect 686 -221 688 -219
rect 690 -221 692 -219
rect 686 -222 692 -221
rect 438 -226 440 -224
rect 442 -226 444 -224
rect 438 -227 444 -226
rect 451 -227 455 -225
rect 451 -229 452 -227
rect 454 -229 455 -227
rect 425 -232 429 -230
rect 425 -234 426 -232
rect 428 -234 429 -232
rect 425 -240 429 -234
rect 451 -232 455 -229
rect 451 -236 475 -232
rect 425 -244 436 -240
rect 432 -250 436 -244
rect 471 -240 475 -236
rect 451 -241 467 -240
rect 451 -243 463 -241
rect 465 -243 467 -241
rect 451 -244 467 -243
rect 471 -242 476 -240
rect 471 -244 473 -242
rect 475 -244 476 -242
rect 451 -250 455 -244
rect 471 -246 476 -244
rect 471 -248 475 -246
rect 432 -251 455 -250
rect 432 -253 434 -251
rect 436 -253 455 -251
rect 432 -254 455 -253
rect 443 -265 447 -263
rect 443 -267 444 -265
rect 446 -267 447 -265
rect 443 -272 447 -267
rect 451 -265 455 -254
rect 459 -251 475 -248
rect 459 -253 460 -251
rect 462 -252 475 -251
rect 462 -253 463 -252
rect 459 -258 463 -253
rect 459 -260 460 -258
rect 462 -260 463 -258
rect 459 -262 463 -260
rect 499 -225 503 -223
rect 508 -224 533 -223
rect 617 -224 642 -223
rect 508 -226 510 -224
rect 512 -225 533 -224
rect 512 -226 530 -225
rect 508 -227 530 -226
rect 532 -227 533 -225
rect 509 -232 524 -231
rect 509 -233 520 -232
rect 495 -234 520 -233
rect 522 -234 524 -232
rect 495 -236 497 -234
rect 499 -235 524 -234
rect 529 -232 533 -227
rect 538 -225 548 -224
rect 538 -227 540 -225
rect 542 -227 548 -225
rect 538 -228 548 -227
rect 529 -234 530 -232
rect 532 -234 533 -232
rect 499 -236 513 -235
rect 529 -236 533 -234
rect 495 -237 513 -236
rect 502 -244 506 -242
rect 502 -246 503 -244
rect 505 -246 506 -244
rect 502 -256 506 -246
rect 509 -248 513 -237
rect 544 -232 548 -228
rect 544 -236 564 -232
rect 560 -239 564 -236
rect 552 -241 556 -239
rect 552 -243 553 -241
rect 555 -243 556 -241
rect 552 -248 556 -243
rect 560 -241 566 -239
rect 560 -243 563 -241
rect 565 -243 566 -241
rect 560 -245 566 -243
rect 509 -252 516 -248
rect 512 -253 516 -252
rect 512 -255 513 -253
rect 515 -255 516 -253
rect 502 -260 508 -256
rect 512 -257 516 -255
rect 560 -256 564 -245
rect 524 -257 564 -256
rect 524 -259 548 -257
rect 550 -259 564 -257
rect 524 -260 564 -259
rect 504 -264 528 -260
rect 547 -264 551 -260
rect 602 -225 612 -224
rect 602 -227 608 -225
rect 610 -227 612 -225
rect 602 -228 612 -227
rect 617 -225 638 -224
rect 617 -227 618 -225
rect 620 -226 638 -225
rect 640 -226 642 -224
rect 647 -225 651 -223
rect 620 -227 642 -226
rect 602 -232 606 -228
rect 586 -236 606 -232
rect 586 -239 590 -236
rect 584 -241 590 -239
rect 584 -243 585 -241
rect 587 -243 590 -241
rect 584 -245 590 -243
rect 586 -256 590 -245
rect 594 -241 598 -239
rect 617 -232 621 -227
rect 710 -226 716 -225
rect 710 -228 712 -226
rect 714 -228 716 -226
rect 710 -229 716 -228
rect 720 -226 726 -218
rect 720 -228 722 -226
rect 724 -228 726 -226
rect 737 -224 752 -223
rect 737 -226 739 -224
rect 741 -226 752 -224
rect 737 -227 752 -226
rect 720 -229 726 -228
rect 617 -234 618 -232
rect 620 -234 621 -232
rect 617 -236 621 -234
rect 626 -232 641 -231
rect 626 -234 628 -232
rect 630 -233 641 -232
rect 630 -234 655 -233
rect 626 -235 651 -234
rect 637 -236 651 -235
rect 653 -236 655 -234
rect 637 -237 655 -236
rect 594 -243 595 -241
rect 597 -243 598 -241
rect 594 -248 598 -243
rect 637 -248 641 -237
rect 634 -252 641 -248
rect 644 -244 648 -242
rect 644 -246 645 -244
rect 647 -246 648 -244
rect 634 -253 638 -252
rect 634 -255 635 -253
rect 637 -255 638 -253
rect 586 -257 626 -256
rect 634 -257 638 -255
rect 644 -256 648 -246
rect 677 -232 695 -231
rect 677 -234 679 -232
rect 681 -234 695 -232
rect 677 -235 695 -234
rect 691 -241 695 -235
rect 691 -243 692 -241
rect 694 -243 695 -241
rect 670 -248 676 -247
rect 586 -259 600 -257
rect 602 -259 626 -257
rect 586 -260 626 -259
rect 642 -260 648 -256
rect 599 -264 603 -260
rect 622 -264 646 -260
rect 691 -256 695 -243
rect 680 -260 695 -256
rect 680 -264 684 -260
rect 698 -264 699 -253
rect 710 -249 714 -229
rect 748 -232 752 -227
rect 755 -224 759 -218
rect 755 -226 756 -224
rect 758 -226 759 -224
rect 755 -228 759 -226
rect 734 -235 745 -233
rect 734 -237 742 -235
rect 744 -237 745 -235
rect 748 -234 762 -232
rect 748 -236 763 -234
rect 734 -239 745 -237
rect 758 -238 760 -236
rect 762 -238 763 -236
rect 734 -249 738 -239
rect 758 -240 763 -238
rect 710 -250 738 -249
rect 710 -252 712 -250
rect 714 -251 738 -250
rect 714 -252 735 -251
rect 710 -253 735 -252
rect 737 -253 738 -251
rect 754 -250 755 -244
rect 734 -255 738 -253
rect 534 -265 540 -264
rect 451 -266 484 -265
rect 451 -268 480 -266
rect 482 -268 484 -266
rect 451 -269 484 -268
rect 534 -267 536 -265
rect 538 -267 540 -265
rect 443 -274 444 -272
rect 446 -274 447 -272
rect 499 -272 505 -271
rect 499 -274 501 -272
rect 503 -274 505 -272
rect 534 -272 540 -267
rect 547 -266 548 -264
rect 550 -266 551 -264
rect 547 -268 551 -266
rect 556 -265 562 -264
rect 556 -267 558 -265
rect 560 -267 562 -265
rect 534 -274 536 -272
rect 538 -274 540 -272
rect 556 -272 562 -267
rect 556 -274 558 -272
rect 560 -274 562 -272
rect 588 -265 594 -264
rect 588 -267 590 -265
rect 592 -267 594 -265
rect 588 -272 594 -267
rect 599 -266 600 -264
rect 602 -266 603 -264
rect 599 -268 603 -266
rect 610 -265 616 -264
rect 610 -267 612 -265
rect 614 -267 616 -265
rect 588 -274 590 -272
rect 592 -274 594 -272
rect 610 -272 616 -267
rect 667 -265 684 -264
rect 667 -267 669 -265
rect 671 -267 684 -265
rect 667 -268 684 -267
rect 758 -257 762 -240
rect 746 -261 762 -257
rect 774 -226 780 -225
rect 774 -228 776 -226
rect 778 -228 780 -226
rect 774 -229 780 -228
rect 784 -226 790 -218
rect 784 -228 786 -226
rect 788 -228 790 -226
rect 801 -224 816 -223
rect 801 -226 803 -224
rect 805 -226 816 -224
rect 801 -227 816 -226
rect 784 -229 790 -228
rect 774 -249 778 -229
rect 812 -232 816 -227
rect 819 -224 823 -218
rect 819 -226 820 -224
rect 822 -226 823 -224
rect 819 -228 823 -226
rect 798 -235 809 -233
rect 798 -237 806 -235
rect 808 -237 809 -235
rect 812 -234 826 -232
rect 812 -236 827 -234
rect 798 -239 809 -237
rect 822 -238 824 -236
rect 826 -238 827 -236
rect 798 -249 802 -239
rect 822 -240 827 -238
rect 774 -250 802 -249
rect 774 -252 776 -250
rect 778 -251 802 -250
rect 778 -252 799 -251
rect 774 -253 799 -252
rect 801 -253 802 -251
rect 818 -250 819 -244
rect 798 -255 802 -253
rect 737 -262 750 -261
rect 737 -264 739 -262
rect 741 -264 750 -262
rect 737 -265 750 -264
rect 822 -257 826 -240
rect 810 -261 826 -257
rect 801 -262 814 -261
rect 801 -264 803 -262
rect 805 -264 814 -262
rect 801 -265 814 -264
rect 610 -274 612 -272
rect 614 -274 616 -272
rect 645 -272 651 -271
rect 645 -274 647 -272
rect 649 -274 651 -272
rect 686 -272 692 -271
rect 686 -274 688 -272
rect 690 -274 692 -272
rect 721 -272 725 -270
rect 721 -274 722 -272
rect 724 -274 725 -272
rect 754 -272 760 -271
rect 754 -274 756 -272
rect 758 -274 760 -272
rect 785 -272 789 -270
rect 785 -274 786 -272
rect 788 -274 789 -272
rect 818 -272 824 -271
rect 818 -274 820 -272
rect 822 -274 824 -272
<< via1 >>
rect 26 291 28 293
rect 159 291 161 293
rect 399 291 401 293
rect 584 291 586 293
rect 776 291 778 293
rect 7 264 9 266
rect 15 244 17 246
rect 47 270 49 272
rect 39 258 41 260
rect 55 247 57 249
rect 79 253 81 255
rect 119 261 121 263
rect 137 253 139 255
rect 87 245 89 247
rect 168 253 170 255
rect 178 266 180 268
rect 208 261 210 263
rect 209 245 211 247
rect 266 270 268 272
rect 257 242 259 244
rect 266 253 268 255
rect 314 270 316 272
rect 298 249 300 251
rect 322 247 324 249
rect 346 253 348 255
rect 386 261 388 263
rect 404 253 406 255
rect 354 245 356 247
rect 435 253 437 255
rect 445 266 447 268
rect 475 261 477 263
rect 476 245 478 247
rect 533 270 535 272
rect 524 243 526 245
rect 533 253 535 255
rect 581 270 583 272
rect 565 249 567 251
rect 589 247 591 249
rect 613 253 615 255
rect 653 261 655 263
rect 671 253 673 255
rect 621 245 623 247
rect 702 253 704 255
rect 712 266 714 268
rect 742 261 744 263
rect 743 245 745 247
rect 800 270 802 272
rect 791 243 793 245
rect 800 253 802 255
rect 832 249 834 251
rect 214 224 216 226
rect 481 224 483 226
rect 748 224 750 226
rect 769 221 771 223
rect 15 193 17 195
rect 55 195 57 197
rect 7 172 9 174
rect 39 181 41 183
rect 79 189 81 191
rect 47 173 49 175
rect 87 197 89 199
rect 137 189 139 191
rect 168 189 170 191
rect 132 181 134 183
rect 259 205 261 207
rect 209 197 211 199
rect 178 176 180 178
rect 226 184 228 186
rect 266 195 268 197
rect 266 176 268 178
rect 322 196 324 198
rect 346 189 348 191
rect 314 173 316 175
rect 290 165 292 167
rect 354 197 356 199
rect 404 189 406 191
rect 435 189 437 191
rect 399 181 401 183
rect 526 205 528 207
rect 476 197 478 199
rect 445 176 447 178
rect 493 184 495 186
rect 533 195 535 197
rect 533 176 535 178
rect 588 194 590 196
rect 613 189 615 191
rect 581 173 583 175
rect 557 165 559 167
rect 621 197 623 199
rect 671 189 673 191
rect 702 189 704 191
rect 666 181 668 183
rect 793 206 795 208
rect 743 197 745 199
rect 712 176 714 178
rect 760 184 762 186
rect 800 195 802 197
rect 800 176 802 178
rect 824 165 826 167
rect 833 147 835 149
rect 8 143 10 145
rect 7 120 9 122
rect 39 117 41 119
rect 47 126 49 128
rect 14 101 16 103
rect 55 104 57 106
rect 79 109 81 111
rect 136 117 138 119
rect 138 109 140 111
rect 87 101 89 103
rect 168 109 170 111
rect 178 122 180 124
rect 226 117 228 119
rect 209 101 211 103
rect 266 126 268 128
rect 266 109 268 111
rect 314 122 316 124
rect 298 105 300 107
rect 322 104 324 106
rect 346 109 348 111
rect 259 93 261 95
rect 403 117 405 119
rect 405 109 407 111
rect 354 101 356 103
rect 435 109 437 111
rect 445 122 447 124
rect 493 117 495 119
rect 476 101 478 103
rect 533 126 535 128
rect 533 109 535 111
rect 581 126 583 128
rect 565 105 567 107
rect 589 104 591 106
rect 613 109 615 111
rect 526 93 528 95
rect 670 117 672 119
rect 672 109 674 111
rect 621 101 623 103
rect 702 109 704 111
rect 712 122 714 124
rect 760 117 762 119
rect 743 101 745 103
rect 800 126 802 128
rect 800 109 802 111
rect 832 105 834 107
rect 793 93 795 95
rect 763 77 765 79
rect 131 74 133 76
rect 14 53 16 55
rect 7 33 9 35
rect 55 54 57 56
rect 39 40 41 42
rect 47 36 49 38
rect 79 45 81 47
rect 87 53 89 55
rect 137 45 139 47
rect 168 45 170 47
rect 131 37 133 39
rect 259 61 261 63
rect 209 53 211 55
rect 178 32 180 34
rect 226 40 228 42
rect 266 51 268 53
rect 266 32 268 34
rect 322 50 324 52
rect 314 32 316 34
rect 346 45 348 47
rect 298 21 300 23
rect 354 53 356 55
rect 404 45 406 47
rect 435 45 437 47
rect 398 37 400 39
rect 526 61 528 63
rect 476 53 478 55
rect 445 32 447 34
rect 493 40 495 42
rect 533 51 535 53
rect 533 32 535 34
rect 589 51 591 53
rect 581 32 583 34
rect 613 45 615 47
rect 565 20 567 22
rect 621 53 623 55
rect 671 45 673 47
rect 702 45 704 47
rect 665 37 667 39
rect 793 61 795 63
rect 743 53 745 55
rect 712 32 714 34
rect 760 40 762 42
rect 800 51 802 53
rect 800 32 802 34
rect 824 21 826 23
rect 25 6 27 8
rect 832 3 834 5
rect 432 -10 434 -8
rect 700 -11 702 -9
rect 441 -37 443 -35
rect 481 -27 483 -25
rect 520 -27 522 -25
rect 540 -35 542 -33
rect 489 -43 491 -41
rect 570 -35 572 -33
rect 580 -22 582 -20
rect 628 -30 630 -28
rect 611 -43 613 -41
rect 668 -22 670 -20
rect 720 -19 722 -17
rect 668 -41 670 -39
rect 719 -43 721 -41
rect 747 -27 749 -25
rect 661 -51 663 -49
rect 776 -19 778 -17
rect 767 -52 769 -50
rect 790 -38 792 -36
rect 806 -27 808 -25
rect 831 -19 833 -17
rect 762 -67 764 -65
rect 436 -91 438 -89
rect 425 -121 427 -119
rect 481 -107 483 -105
rect 489 -91 491 -89
rect 539 -99 541 -97
rect 570 -99 572 -97
rect 526 -107 528 -105
rect 661 -83 663 -81
rect 611 -91 613 -89
rect 580 -112 582 -110
rect 628 -107 630 -105
rect 668 -99 670 -97
rect 700 -95 702 -93
rect 668 -116 670 -114
rect 718 -91 720 -89
rect 767 -91 769 -89
rect 750 -107 752 -105
rect 719 -115 721 -113
rect 806 -107 808 -105
rect 775 -115 777 -113
rect 831 -110 833 -108
rect 835 -142 837 -140
rect 426 -161 428 -159
rect 481 -171 483 -169
rect 434 -188 436 -186
rect 521 -171 523 -169
rect 540 -179 542 -177
rect 489 -187 491 -185
rect 570 -179 572 -177
rect 580 -166 582 -164
rect 628 -174 630 -172
rect 611 -187 613 -185
rect 668 -166 670 -164
rect 718 -163 720 -161
rect 668 -185 670 -183
rect 700 -184 702 -182
rect 718 -187 720 -185
rect 745 -171 747 -169
rect 776 -163 778 -161
rect 767 -171 769 -169
rect 661 -195 663 -193
rect 807 -172 809 -170
rect 831 -170 833 -168
rect 765 -211 767 -209
rect 435 -234 437 -232
rect 426 -257 428 -255
rect 481 -251 483 -249
rect 489 -235 491 -233
rect 540 -243 542 -241
rect 570 -243 572 -241
rect 531 -251 533 -249
rect 661 -227 663 -225
rect 611 -235 613 -233
rect 580 -256 582 -254
rect 622 -251 624 -249
rect 668 -243 670 -241
rect 668 -256 670 -254
rect 700 -239 702 -237
rect 718 -235 720 -233
rect 749 -251 751 -249
rect 814 -251 816 -249
rect 767 -255 769 -253
rect 712 -268 714 -266
rect 831 -251 833 -249
rect 776 -268 778 -266
rect 461 -282 463 -280
rect 529 -281 531 -279
rect 612 -281 614 -279
rect 709 -281 711 -279
rect 773 -281 775 -279
<< via2 >>
rect 31 292 33 294
rect 164 292 166 294
rect 404 292 406 294
rect 589 292 591 294
rect 781 292 783 294
rect 53 270 55 272
rect 305 270 307 272
rect 574 270 576 272
rect 1 264 3 266
rect 211 261 213 263
rect 333 261 335 263
rect 478 261 480 263
rect 600 261 602 263
rect 745 261 747 263
rect 43 247 45 249
rect 302 249 304 251
rect 21 244 23 246
rect 310 247 312 249
rect 569 249 571 251
rect 577 247 579 249
rect 836 249 838 251
rect 262 242 264 244
rect 529 243 531 245
rect 755 243 757 245
rect 211 224 213 226
rect 478 224 480 226
rect 745 224 747 226
rect 773 221 775 223
rect 333 205 335 207
rect 600 205 602 207
rect 789 206 791 208
rect 1 193 3 195
rect 62 195 64 197
rect 290 196 292 198
rect 555 194 557 196
rect 302 184 304 186
rect 569 184 571 186
rect 836 184 838 186
rect 321 181 323 183
rect 589 181 591 183
rect 15 172 17 174
rect 43 173 45 175
rect 310 173 312 175
rect 577 173 579 175
rect -9 133 -7 135
rect 64 126 66 128
rect 1 120 3 122
rect 299 122 301 124
rect 568 126 570 128
rect 834 152 836 154
rect 334 117 336 119
rect 600 117 602 119
rect 43 104 45 106
rect 302 105 304 107
rect 310 104 312 106
rect 569 105 571 107
rect 577 104 579 106
rect 836 105 838 107
rect 23 101 25 103
rect 321 93 323 95
rect 589 93 591 95
rect 801 93 803 95
rect 767 77 769 79
rect 127 74 129 76
rect 334 61 336 63
rect 601 62 603 64
rect 811 61 813 63
rect 31 53 33 55
rect 62 54 64 56
rect 43 48 45 50
rect 290 50 292 52
rect 552 51 554 53
rect 1 33 3 35
rect 302 40 304 42
rect 569 40 571 42
rect 836 40 838 42
rect 127 37 129 39
rect 394 37 396 39
rect 661 37 663 39
rect 310 32 312 34
rect 577 32 579 34
rect 39 20 41 22
rect 394 21 396 23
rect 661 20 663 22
rect 821 21 823 23
rect 20 6 22 8
rect 833 8 835 10
rect 39 2 41 4
rect 405 2 407 4
rect 390 -10 392 -8
rect 577 -10 579 -8
rect 541 -29 543 -27
rect 704 -30 706 -28
rect 730 -19 732 -17
rect 831 -22 833 -20
rect 751 -27 753 -25
rect 789 -28 791 -26
rect 418 -37 420 -35
rect 767 -46 769 -44
rect 766 -67 768 -65
rect 418 -91 420 -89
rect 704 -95 706 -93
rect 767 -95 769 -93
rect 490 -99 492 -97
rect 692 -107 694 -105
rect 745 -107 747 -105
rect 801 -107 803 -105
rect 730 -115 732 -113
rect 831 -114 833 -112
rect 310 -121 312 -119
rect 529 -128 531 -126
rect 744 -128 746 -126
rect 835 -139 837 -137
rect 262 -150 264 -148
rect 748 -150 750 -148
rect 51 -161 53 -159
rect 730 -163 732 -161
rect 831 -167 833 -165
rect 748 -171 750 -169
rect 704 -174 706 -172
rect 767 -174 769 -172
rect 811 -172 813 -170
rect 508 -179 510 -177
rect 418 -188 420 -186
rect 692 -184 694 -182
rect 769 -211 771 -209
rect 418 -234 420 -232
rect 704 -239 706 -237
rect 464 -243 466 -241
rect 618 -251 620 -249
rect 746 -251 748 -249
rect 767 -251 769 -249
rect 821 -251 823 -249
rect 1 -257 3 -255
rect 831 -255 833 -253
rect 730 -268 732 -266
rect 418 -271 420 -269
rect 618 -271 620 -269
rect 466 -282 468 -280
rect 534 -282 536 -280
rect 617 -282 619 -280
rect 714 -282 716 -280
rect 778 -282 780 -280
<< via3 >>
rect 31 303 33 305
rect 164 303 166 305
rect 404 303 406 305
rect 589 303 591 305
rect 781 303 783 305
rect 31 283 33 285
rect 21 221 23 223
rect -9 136 -7 138
rect 15 149 17 151
rect 23 77 25 79
rect 53 283 55 285
rect 305 283 307 285
rect 464 283 466 285
rect 62 221 64 223
rect 64 149 66 151
rect 62 77 64 79
rect 20 9 22 11
rect 1 -51 3 -49
rect 51 -41 53 -39
rect 290 221 292 223
rect 299 149 301 151
rect 290 77 292 79
rect 390 -14 392 -12
rect 310 -28 312 -26
rect 405 -260 407 -258
rect 574 283 576 285
rect 508 221 510 223
rect 490 149 492 151
rect 555 221 557 223
rect 568 149 570 151
rect 541 77 543 79
rect 552 77 554 79
rect 777 221 779 223
rect 771 77 773 79
rect 845 152 847 154
rect 767 -42 769 -40
rect 770 -67 772 -65
rect 767 -99 769 -97
rect 767 -177 769 -175
rect 773 -211 775 -209
rect 767 -247 769 -245
rect 844 8 846 10
rect 862 -1 864 1
rect 831 -25 833 -23
rect 831 -118 833 -116
rect 846 -139 848 -137
rect 831 -164 833 -162
rect 746 -260 748 -258
rect 831 -259 833 -257
rect 870 -9 872 -7
rect 878 -17 880 -15
rect 878 -118 880 -116
rect 870 -164 872 -162
rect 862 -259 864 -257
rect 730 -273 732 -271
rect 466 -293 468 -291
rect 534 -293 536 -291
rect 617 -293 619 -291
rect 714 -293 716 -291
rect 778 -293 780 -291
<< via4 >>
rect 28 303 30 305
rect 161 303 163 305
rect 401 303 403 305
rect 586 303 588 305
rect 778 303 780 305
rect 782 221 784 223
rect 845 149 847 151
rect -9 139 -7 141
rect 775 77 777 79
rect -9 9 -7 11
rect 844 5 846 7
rect 774 -67 776 -65
rect 846 -143 848 -141
rect 778 -211 780 -209
rect 463 -293 465 -291
rect 531 -293 533 -291
rect 614 -293 616 -291
rect 711 -293 713 -291
rect 775 -293 777 -291
<< via5 >>
rect 810 220 814 224
rect 810 76 814 80
rect 809 -68 813 -64
rect 809 -212 813 -208
<< labels >>
rlabel alu1 214 226 214 226 1 gnd
rlabel alu1 214 218 214 218 5 gnd
rlabel alu1 132 218 132 218 5 gnd
rlabel alu1 237 290 237 290 1 Vdd
rlabel alu1 263 290 263 290 1 Vdd
rlabel alu1 173 290 173 290 1 Vdd
rlabel alu1 108 290 108 290 1 vdd
rlabel alu1 108 153 108 153 1 Vdd
rlabel alu1 173 154 173 154 1 Vdd
rlabel alu1 264 154 264 154 1 Vdd
rlabel alu1 238 154 238 154 1 Vdd
rlabel alu1 238 10 238 10 1 Vdd
rlabel alu1 264 10 264 10 1 Vdd
rlabel alu1 173 10 173 10 1 Vdd
rlabel alu1 108 9 108 9 1 Vdd
rlabel alu1 108 146 108 146 1 vdd
rlabel alu1 173 146 173 146 1 Vdd
rlabel alu1 263 146 263 146 1 Vdd
rlabel alu1 237 146 237 146 1 Vdd
rlabel alu1 132 74 132 74 5 gnd
rlabel alu1 214 74 214 74 5 gnd
rlabel alu1 214 82 214 82 1 gnd
rlabel alu1 132 82 132 82 1 gnd
rlabel alu1 64 146 64 146 4 vdd
rlabel alu1 64 154 64 154 2 vdd
rlabel alu1 24 154 24 154 2 vdd
rlabel alu1 24 290 24 290 4 vdd
rlabel alu1 8 270 8 270 1 b_0
rlabel alu1 48 175 48 175 1 b_1
rlabel alu1 8 179 8 179 1 a_2
rlabel via1 16 194 16 194 1 b_0
rlabel alu1 16 248 16 248 1 a_1
rlabel alu1 56 194 56 194 1 a_1
rlabel alu1 24 146 24 146 4 vdd
rlabel alu1 8 122 8 122 1 b_0
rlabel alu1 16 105 16 105 1 a_3
rlabel alu1 56 106 56 106 1 b_1
rlabel alu1 48 122 48 122 1 a_2
rlabel alu1 8 33 8 33 1 b_0
rlabel alu1 16 50 16 50 1 a_0
rlabel alu1 40 45 40 45 1 p_0
rlabel alu1 56 50 56 50 1 a_3
rlabel alu1 48 34 48 34 1 b_1
rlabel alu1 48 266 48 266 1 a_0
rlabel alu1 258 259 258 259 1 p_1
rlabel alu1 481 226 481 226 1 gnd
rlabel alu1 481 218 481 218 5 gnd
rlabel alu1 399 218 399 218 5 gnd
rlabel alu1 504 290 504 290 1 Vdd
rlabel alu1 530 290 530 290 1 Vdd
rlabel alu1 440 290 440 290 1 Vdd
rlabel alu1 375 290 375 290 1 vdd
rlabel alu1 375 153 375 153 1 Vdd
rlabel alu1 440 154 440 154 1 Vdd
rlabel alu1 531 154 531 154 1 Vdd
rlabel alu1 505 154 505 154 1 Vdd
rlabel alu1 505 10 505 10 1 Vdd
rlabel alu1 531 10 531 10 1 Vdd
rlabel alu1 440 10 440 10 1 Vdd
rlabel alu1 375 9 375 9 1 Vdd
rlabel alu1 375 146 375 146 1 vdd
rlabel alu1 440 146 440 146 1 Vdd
rlabel alu1 530 146 530 146 1 Vdd
rlabel alu1 504 146 504 146 1 Vdd
rlabel alu1 399 74 399 74 5 gnd
rlabel alu1 481 74 481 74 5 gnd
rlabel alu1 481 82 481 82 1 gnd
rlabel alu1 399 82 399 82 1 gnd
rlabel alu1 331 146 331 146 4 vdd
rlabel alu1 331 154 331 154 2 vdd
rlabel alu1 323 194 323 194 1 a_1
rlabel alu1 315 122 315 122 1 a_2
rlabel alu1 323 50 323 50 1 a_3
rlabel alu1 315 266 315 266 1 a_0
rlabel via1 323 248 323 248 1 b_2
rlabel via1 315 175 315 175 1 b_2
rlabel via1 323 106 323 106 1 b_2
rlabel via1 315 34 315 34 1 b_2
rlabel alu1 748 226 748 226 1 gnd
rlabel alu1 748 218 748 218 5 gnd
rlabel alu1 666 218 666 218 5 gnd
rlabel alu1 771 290 771 290 1 Vdd
rlabel alu1 797 290 797 290 1 Vdd
rlabel alu1 707 290 707 290 1 Vdd
rlabel alu1 642 290 642 290 1 vdd
rlabel alu1 642 153 642 153 1 Vdd
rlabel alu1 707 154 707 154 1 Vdd
rlabel alu1 798 154 798 154 1 Vdd
rlabel alu1 772 154 772 154 1 Vdd
rlabel alu1 772 10 772 10 1 Vdd
rlabel alu1 707 10 707 10 1 Vdd
rlabel alu1 642 9 642 9 1 Vdd
rlabel alu1 642 146 642 146 1 vdd
rlabel alu1 707 146 707 146 1 Vdd
rlabel alu1 797 146 797 146 1 Vdd
rlabel alu1 771 146 771 146 1 Vdd
rlabel alu1 666 74 666 74 5 gnd
rlabel alu1 748 74 748 74 5 gnd
rlabel alu1 748 82 748 82 1 gnd
rlabel alu1 666 82 666 82 1 gnd
rlabel alu1 598 146 598 146 4 vdd
rlabel alu1 598 154 598 154 2 vdd
rlabel alu1 590 194 590 194 1 a_1
rlabel alu1 582 122 582 122 1 a_2
rlabel alu1 590 50 590 50 1 a_3
rlabel alu1 582 266 582 266 1 a_0
rlabel via1 590 248 590 248 1 b_3
rlabel via1 582 175 582 175 1 b_3
rlabel via1 590 106 590 106 1 b_3
rlabel via1 582 34 582 34 1 b_3
rlabel alu1 792 46 792 46 1 p_6
rlabel alu1 792 115 792 115 1 p_5
rlabel alu1 792 190 792 190 1 p_4
rlabel alu1 792 259 792 259 1 p_3
rlabel alu1 525 259 525 259 1 p_2
rlabel alu1 798 10 798 10 1 Vdd
rlabel alu1 804 -142 804 -142 4 vdd
rlabel alu1 807 -205 807 -205 1 gnd
rlabel alu1 777 -153 777 -153 1 sel
rlabel alu1 713 -153 713 -153 1 sel
rlabel alu1 743 -205 743 -205 1 gnd
rlabel alu1 740 -142 740 -142 4 vdd
rlabel via1 777 -267 777 -267 5 sel
rlabel alu1 807 -215 807 -215 5 gnd
rlabel alu1 804 -278 804 -278 2 vdd
rlabel alu1 740 -278 740 -278 2 vdd
rlabel alu1 743 -215 743 -215 5 gnd
rlabel via1 713 -267 713 -267 5 sel
rlabel alu1 713 -123 713 -123 5 sel
rlabel alu1 743 -71 743 -71 5 gnd
rlabel alu1 740 -134 740 -134 2 vdd
rlabel alu1 804 -134 804 -134 2 vdd
rlabel alu1 807 -71 807 -71 5 gnd
rlabel alu1 777 -123 777 -123 5 sel
rlabel alu1 740 2 740 2 4 vdd
rlabel alu1 743 -61 743 -61 1 gnd
rlabel alu1 777 -9 777 -9 1 sel
rlabel alu1 807 -61 807 -61 1 gnd
rlabel alu1 804 2 804 2 4 vdd
rlabel alu1 546 -98 546 -98 5 a_2
rlabel alu1 546 -34 546 -34 5 a_3
rlabel alu1 660 -34 660 -34 5 s_3
rlabel alu1 660 -103 660 -103 5 s_2
rlabel alu1 534 -70 534 -70 5 gnd
rlabel alu1 616 -70 616 -70 5 gnd
rlabel alu1 701 -28 701 -28 1 cout
rlabel alu1 616 -62 616 -62 1 gnd
rlabel alu1 534 -62 534 -62 1 gnd
rlabel alu1 639 -134 639 -134 5 Vdd
rlabel alu1 665 -134 665 -134 5 Vdd
rlabel alu1 575 -134 575 -134 5 Vdd
rlabel alu1 510 -134 510 -134 5 vdd
rlabel alu1 510 3 510 3 5 Vdd
rlabel alu1 575 2 575 2 5 Vdd
rlabel alu1 666 2 666 2 5 Vdd
rlabel alu1 640 2 640 2 5 Vdd
rlabel alu1 640 -142 640 -142 5 Vdd
rlabel alu1 666 -142 666 -142 5 Vdd
rlabel alu1 575 -142 575 -142 5 Vdd
rlabel alu1 510 -141 510 -141 5 Vdd
rlabel alu1 510 -278 510 -278 5 vdd
rlabel alu1 575 -278 575 -278 5 Vdd
rlabel alu1 665 -278 665 -278 5 Vdd
rlabel alu1 639 -278 639 -278 5 Vdd
rlabel alu1 660 -247 660 -247 5 s_0
rlabel alu1 660 -178 660 -178 5 s_1
rlabel alu1 546 -178 546 -178 5 a_1
rlabel alu1 546 -242 546 -242 5 a_0
rlabel alu1 534 -206 534 -206 1 gnd
rlabel alu1 616 -206 616 -206 1 gnd
rlabel alu1 613 -250 613 -250 5 cin
rlabel alu1 616 -214 616 -214 5 gnd
rlabel alu1 534 -214 534 -214 5 gnd
rlabel alu1 832 -34 832 -34 1 out_4
rlabel alu1 832 -104 832 -104 1 out_5
rlabel alu1 833 -174 833 -174 1 out_6
rlabel alu1 831 -248 831 -248 1 out_7
rlabel alu1 768 -31 768 -31 1 out_3
rlabel alu1 454 2 454 2 6 vdd
rlabel alu1 454 -134 454 -134 8 vdd
rlabel alu1 454 -142 454 -142 6 vdd
rlabel alu1 454 -278 454 -278 8 vdd
rlabel alu1 426 -18 426 -18 1 b_3
rlabel alu1 426 -114 426 -114 1 b_2
rlabel polyct1 442 -38 442 -38 1 cin
rlabel alu2 434 -90 434 -90 1 cin
rlabel via1 434 -186 434 -186 1 cin
rlabel alu2 434 -234 434 -234 1 cin
rlabel alu1 768 -101 768 -101 1 out_2
rlabel alu1 433 -266 433 -266 1 b_0
rlabel alu1 57 252 57 252 1 b_1
rlabel alu1 426 -164 426 -164 1 b_1
rlabel alu1 833 48 833 48 1 p_7
rlabel alu1 764 -154 764 -154 1 out_1
rlabel alu1 769 -196 769 -196 1 out_1
rlabel alu4 -42 -272 -42 -272 1 sel
rlabel alu1 769 -224 769 -224 1 out_0
rlabel alu1 769 -261 769 -261 1 out_0
rlabel alu1 716 -18 716 -18 1 sel
rlabel alu4 -48 224 -48 224 1 a_1
rlabel alu4 -47 199 -47 199 1 a_3
rlabel alu4 -47 211 -47 211 1 a_2
rlabel alu4 -48 233 -48 233 1 a_0
rlabel alu4 -71 -50 -71 -50 3 b_0
rlabel alu4 -71 -40 -71 -40 3 b_1
rlabel alu4 -70 -27 -70 -27 3 b_2
rlabel alu4 -70 -13 -70 -13 3 b_3
rlabel alu4 901 -24 901 -24 1 out_4
rlabel alu4 903 -16 903 -16 7 out_5
rlabel alu4 901 -8 901 -8 1 out_6
rlabel alu4 901 -1 901 -1 1 out_7
rlabel alu4 901 -41 901 -41 1 out_3
rlabel alu4 902 -49 902 -49 1 out_2
rlabel alu4 903 -58 903 -58 7 out_1
rlabel alu4 903 -65 903 -65 7 out_0
<< end >>
